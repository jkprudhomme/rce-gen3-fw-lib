XlxV64EB    fa00    1f50���r<s1=I%ĨEĿ��|���t�������d\�s��a�#J�N��|��	G�>;��n��&�6���@��)�P�Ֆ�B��`-�Tfh	��6J��h��O�*.�d[Z��<��)�H��UK���J�����;ٍ�����i瞦�
l.*���j?��=F�I�{���Ń�����mmV��@'�q��P��J�������L�l�֓�}d�擖��5�f�q�6���ԓw�X����N��Dﰾ�y��\!���s{Q��XR�=x��UW�x�5ힲv�SR����}������Q�C�Q�3_��W���sE8��y�@ف������ظW������-$w��.f�-*yK�k�ܓ1B=~3�&��,���1�(��Y�����}oܵ��V�cV�������}M)�-14G�)A\+w!��=����U +{��i������v��R�Q��P'k�ߴ�FW�rfq��<�G�|��JM]zT��v���3�s�ɳ�Kd5QAU�Z��6���H��O�Tv����hN�b�/�/����A���^&�\.�p������\��1���8��3��}��r�TW��u�'Ҏ+ɜ�Ҵ)��2�����o�3$�
0� 0)�)�C�K@;��+Q/�U\�r���<�A���*F*�>SxZ=H&�΋"� ��'�
E���Vn�qf�5���t�<u�ʲ��g�^״({N�gh ��{�ӂ�Sy^Q���j�Y�5�@�Ya��sW>�Ah��W��|�6����"�fq�4�U��{�.�#l��ބ�5;G��o�e�GS��WJ�,A*�\�M���2p�o�gW�	�N��6T/�s�	�{��W���_�@�Xr�^���44�� mi��ܦ���ws5ѳP�媝g+���%Yw��1�uoZsq����M���ŀd��Iv1�j_�v�|.����xiu6p/h�,����8�س<���U�X��G�U�Ū�u|��XAe�>^ZlE�ա�2bz�r���OCZ~-��t��(-M�`W���5� d��)ömXl�K��K�	@j[xj���/��e��ġ�-�@�1�Q�>�.r����2T�3��J�e�-�}�M��5N[|\�	�#JJ�wY��2c��m4�O/\ ]�u�[I�@�XW���z���M�����z2�AԹ��li��AB�VV��ҥ��}%+v�lP���|	֪�17{�~�(�&�����96ˑŁ���DNҊLfk� �����#s1!��{'���0X����CE����
:�6����@�3)�4�`���1�#������>�
��ULJԉ��|E����CN�w�E�<�OF����ө�f�c"ӣ�"�@^�.�"��}�#p>o床46Sr��W��G��Y�*��u�q�a��^��RΊ�j��?�)K�'`�75'�V�Oz��=���y�x�+�hz��d��KϜ�h���\��ńS^���bx[Ͼg���t垔P-
��"����6�,;:@k�A��71�ik�MI��>s�1:8p�6��h��|p��5M!p߱��'�T��*nZ��ܝ X�X�����T��cņ��H�o~����A�j�jP��X�?��x-^S���H�^���eC�ُ���	� ;����ߗ^��tv:�gŸ���\�ḵ�F=1�+P_�TfAh�T�W{��.�{�Wl�@��Ҕ��z�'�ɷ~�? �Z�42�F�^m���҄�$$�7+��@��+
�L0'�I���Aξ��I��c?>�PIA\o�:*I�c���|��5�@MP���0iF/�`�;�̇�iK�6SV�w�B���	� �U�*L��� �KB4	I��/Ș�N�+v��R�ܤ��D�6��)���r8��i4��v� ��:n�'f�������wm6?��?7�����-��j��`S�
ў"�o����O��v�(z񉉙�W�;�l(D<���v�`N6��)��4��#k>��FtK��7Q����m/O�x�h��'���7����sHm^��*)�b���m�t��9���Aw�a~e��1X�6��OZ�ʾ��m��[e��p�K��|x}]���XX��1u/_ڿ��%"�8o��Q���T#���٢Z�B������x\+�w�"�~(���.w�l��=k\d��˷R�Z����m�m\��.�pM�92Ƒ^���"�D:=�+=mS��a�rǒ$ֲ�=�]!����
���c�I���g4Z���8  �d
՛�&��i�����2�m8h��A���0)Oq�LX7��U(��b�}l��E�j��~���`<yiy��������|��E�</H�W�£M��lU���[���A�(@�xui�*?��wߏ�E$P�"��Z���eA�u �A�5�~_V�)��Z�>U:)B!������]�=���%y���+�_��_������5)�]_�;�I�M�t��iD�F���D>,�����9�z�g{����w^���y=�gwn�y�P��^4���"$�����C��;<����+ѵ�DV�?�Å��'���߅�3A���d/��Wv%6��O;�����͸����t�ᤂ��B\J�(�x]�e��O΢@�D��<��Ry�ԕ�q����t:1��2���Ӓ�j;�e�6�ySv�ͧoVO�x��7����,��8��`��B�b��1��+�I����KE�����>�\;K��_�v������<^,W1��<s���.�N:kⷁ�r��Pc6�0����^H�
���)�#��L4�Ǥ�������#e�8^�oo
��EŅ�>���E9x�,��^��M�X�=ּ=q�*�d�Mu���Y�� etEy�fǠ�x��sS*Bg���O����+v+	����ת�X���I��5�`�%���)g�]*������%I�ȇ\�����KS�4W6Tj���z��������ը�T/�F���Ѯ�,�R��U�MIA2���$�S�y�K~��x]g'U8��ˤy��7uT�q�xXcw�힬�S��{ k0!��}�}Q�V6B|�mq��Z&���
$�*���+Je�Z�Q:��7�u�A5��i`�ޣM2�C�C~�8M���LҼ�q�e(�(��b������-��I���i�8�=��е����C�q����?+�����Z	fT*���p���A���_:�2t�ze��B���`6'm�|(�'�B+c�Mܵ`'VK?�YX6˘�*��=��)�m�d�8�P�( _)d�c/y��8�LA�]�|�N��i���������`�kxN <(���ӑ���kP�l�;��=��'��$�aQ��ҌZɐKGC�<�87.��t��֬6�;�B�ԩ;`:k#����~Kdy䪍�i�ؽz�r���ˀ��w���W����3�R�l�����*�@�L+F+�<L�r�Z��H�c����yrw��R�h"q\gB�Q��wZY/���Nx�\�gϵzc �Oi�{k�v٦����6"��Px���~��+42[ˋhx��ޑ?L��L}��P82�m��A��g&8���IZ��(����B0Go�Ω��e�.��bl��� 3Q�d�'��B�r#h��lxo�S9?�yDNj��?�ЩM���Ŷ+!���)�Cu��w���[�4��!KSv'\w���P���/dq�4|`�M��󰂜��kN���`v��zKா�Z[.W?R���=g���M��¡�P��oFT��@�}_�[�>���(5�[U�M{[�Ap�X�G��o�Y�4�x@`����]�F�!d�0Dʎg[���d�� !�����ȎB(Zw}���e��]V�IyS�	�l:�.H���s��r����>ߧ��`�j>��@�����X��[Qe�9/6����=� w���Z(�"��> �ud$�����%u�m:%�V����v��[�Z��k�����݋�����[�U��Kc���������v_!�l(����&�ug�6J���?{��J�5V����N�]�:�P�p^���+�; ԯ6�("�ꉣђ�[��M#��o>mq<�#ܡ�<�#��1�����ʗ��C�~R����`���G�X���r��͢|�o��T,P��6м-[���N�	��P���L
m:\�+�kX�EyO�dɦ�Ҩ���;��2��٭��u�V��P�ɣ.#n乨�J�!}�5���))�+�C�}} �I[-�5����J���^}?�����?�b����0Ԃ%���h�h�zڦ�K�ߍ���d�Xz&yB�b�	�(���z����Gp��纻Y폢���L��nc����e+�	�����\�q�B��_<F����<�&nٓR�Jtn��hOb�N#Wj׳�U�����tr֙J�"��8Z�� ���������s&(����+�v�nK���D�ъ�#��?�aǡ����8�j�Lē��8���C��f��k0 ��z�<�S�˥bC��'R<w+�Q�ғ�vqd�j9辌ƈp�����b�ρ����0� ��G%1uמnU"�އ̀��L�Q�]	c|$�m|�`�%�z����]��M��R\xw�����G{��C3 ��P�7�e��k���r�^*�'���D(Q1���Ͱ�9������8z��<���}���D������}Jy"1�B2�1Y<j��},�Rb���L��b*�q|��o ��:LCib��)��auH]�Ⱥ���e��Ǔʮ�*�Dn�#T�,��;}�(�zLO��=�g��Q5BO�Gv��H7��5�N�>�5���X<�-=�t6�;+ �$�������j�KG�ґ�����Ʈ0mI.���Ƃa��ò��p��UˣYR*���{ ��s��0b�\�n_��y�G&�,o�^�=�����r��I#8�e[
NCZ���Go4�}}I�qp9%T��E�(�0����:f���jsa�2wM7��t�sm��P���v�1i��פ�_��/X	Ql2���e�,��WD�x���p7X��C��zO 	L�Ԩ(�����jsVtv�5	��D���#�!e�y���P�	$H��]�,��>P��r,�'��?��-l�:x8� ���M;�J� xMDL\B
�Sڰ�#h�j!�VZ#����3��3
�a�j�5~dK�˒0���aK��(���#&��q_kh�"��.
zx�fK��g*����_��^uyd�%�������3�������KG�y]<�5 wgB�'�yvȥ+��+��rϯ���7O�/Eu�Pk�齾�d}�b�ܥ`oTw�|��M��BsPM��~���-�^4��j:Ç�M3�5���G���譼����O��<n�0�6ւ eC"������v�M��*Q=�\��9e�W��8Ꝋ�n��*�"�2=<��&&24�+Sz=T�>�o������v60$��pw���zwi�ۈhU\�m��Ekc�p03l��[E����
.-��c�
+���zx�r�@=�̗J��G̸�,��� �}y-m�k�"��|��k�]�0Z�6O��Ǆ�_�\�z߼��~�,����t�?A8_�$tz$mfL65��P%��:HM�b�DO���P1s{�+���Ñ�4���W��В���X��p[�D���`�"��Re�Ы�4���}������P"�V�:(X��w1h^)���̸'O%mϝY���	('U�W���I5������鯺�gE<�er�,߄;�F$9��g<�7�,��m��у�TUU�4��v�64�G��&m~���L�3b�i��~10��2]�T�t�~b*�F��7��M�D�ACR�M������o���l�2����_qגp��F9pQ���\�.|_>�ہ�+a�a7V\a��=������$����W��ن[�sKL8t�Q��� Vߊ�3gn���c�}�$Y�4�М�PCͥ��50��RdN���!C�s�9�r=��¡�����M7%?���O,}lǙ|�ީ��A�*N�5���s�s�;=�bh��Q��j��M�~�R~ -
��B��0:G��"P>��w�()���n�>�ń8[���Z�n[��EH����0��w��R���N؝�ߚgSSD;I��D�W��~�&��.����e�OE7H��Ԥ �� �H��h�k&c��
�s6k_u��#�z�s�a�(���g�U�QG�V#�dh蠪�g
g�q3��B�.��%d�?g^0ؘ(�N�ſ���#5��e,��eNm�^\�;ڜzzǏ�qŸ���<�7�=yC�
�=�����"�]����[�Ӏ�Ä(܂<ԋޥ���e����b��*N��Ɋ� [n�����:�%\��KN��6;��r4�L���Tdl(�S�\�o�@H�v# �J˹�hKǨ��nh�!��.J`l�c��<��m��k�G@�O}��Ч3��4차�֒���L �7�DW�F�O�Z�m+�q�/P�ǂ�"��x�)�����׸8Dq"�1]�Na��"MՓ��,��m�(�-��Q''0u�m�|~�éu�ኻ��m����=J���+����線:��H!�ᕂQ\g"=���z�������Ü�z���2l�!`��l5��,���*���:�4�yI�V��w�!�����hi�DCa� �8��֊�m�&�Sa]:V	�rc��]����7l���Ul0�M���D���x^���JZ�Ӊ]�pu�c�?�+�f�e��LZq�ѷ���97�	  ��-���H �řa��J�J�S�:�7���}�\jŕ���Ȟ�a�+���X���Z\�p��˛�}�(f�����ur��E����{�5H+H�f�>VpfZ�cJArWŲ�������x7��^-�!�2��V��-mqBH�E���Y<���z㑠��y�vU��6
k�����,�c�Y��/�6c�q�{^Y���ީHg�Z*uc��b����T~P�yJ�:*�������ރ3Nq��>j��+�u�}s��찹P	b�m7黮A��N0�e�Q]��
B	�=���Cҥ�d���ِ��ܟb���UM6���lV�L��HXj��Z�>��A}�;MV�a�L��dZ���r�59�o�?�tj����-a�^b��P�b��8�f�{[�p��x�W�3f2�T5�р�0�(���Z3���Ƞ�.N��Hp��p�	�}!;8Q`p�"�-V\�8��U�m�Ӂgë����u�J����\+�w��ydC%S!��M�c�(�$�����+ ,t��,��^�BcHh/�|�bt�R�)�&%m�n���E�i��x۸<�ܬ{ܖ�Y����n��C�P�|��F�� ����w��t��D}�i�q+�����OKz��\��LQq���!�'���������-X��!m Ͻ]dF_#w�b�L�s�8v��Q�K��*�L)��˓Ҟ|�炉�"y���mf��T\����q8T�x=�7�KM�tv�l'�G���6�]!v^���v?�;K�v����QM����� ���ܛ�*���ɥ�=Ab���^�F[�l4����F��R(�^�:�d(&R�~r��*ϓ��E�ֽ�+�T�nJ��iА�c��,��	z����>�0�iXg gd9���?HR�df���T�R��%���������֏	��`�/�H%�o(�{Y�CVe V0�`A�����z9����=�O��.�*�ʁ�����`Œ�Υ��|y-�ڗ��������×I�b(��:����f �(�I偀ޑq�%�(;R���\[�x�\d�e��k
IT�>���GW�}i&���(ݩ���!΃�(��aXlxV64EB    3367     810���H������yf/�ޯ�#']B��'���v�џɝ���>����ɤ�яס����]�M�����Ғ��Z�N������T���)�P� ���e2G��:<�9��������z����u)�&x�ź�M�:ß����BW�Z�s����/����Bs�ώ�c��:4'}��[���]�4�5g��6�A貚�O)�g>U�%*Ѳ��ZSҵQ�ҋ��WM3��
�����ƀ
C3Rƈ~��C���킿�SOu�	cp^:
�nP�!�����ϒ�`���{q��4��1����x�Rv=���������z
����aT�HO�!��\KMrهw�J����3�`8C O�Xj��d�ğk�6�f�F�̖�;���	�gL��	��$Ή+r�GFo6���y�R�JA΀����aB}$�b��j���gO{km�X�E�$X7a�[���L>&��X:4����P��[�zh<��\za���1]\QQ���c�L�!;L%;����6{�����V+D2��6��Op��Hڋ�{
�q�VM��N��q���#q���<^�u���B����-�����T�&$|��!�fE a�(f��d��d�bk��V'5�FY��-9��w���>\g����2��+��Vm�$����4j��� ̊���*�ÞS$ĭ���l�_�a9������8x*� ��;�:�H����M������X�p���TV���u�i	�;�҂���G$tD�&�����| 8�%��+S���n}�������rˍ��'74��'���E-8�x�װ���p��Z��_%h�y �&�?8�������O���s#�޺j�=���s`�X�rC0bIJ�q�H�]��>#v�X��
-`����1�լ�[b���������`�*?-L����K$�?�Δ�[�r�P��3��֑I)���;}l�ne<D�	���$��3�����x|��&�a:č@C���n�c�C�X_*������o���<l���~�����l�u�	3�+|jn��b��i�8�E#3*�w�� �5�`E(�l����	"���V�%	��o��6'�������kq��^�=�,�@y�r8�;b9 ����e����}oc�!�*�d�_�5��0'��Jq�ڥ1�<s���~��G~M�9�M}�%x��U��b�q.�Zފ�G�PAYᘅ��~�?������-Ʋd���d|T����Ώ%7{�e�U�$Em#'[^%^I]� k%���$M� �bt��\��%�?}O;��(�{�� �5GȪ��}�i̡M��=c!	�k!\�~;�b�h$��O	�X8�`}B�N�@_j�yt�°���,3,k#����B�3`o�hr�#�#��i�3��R3��S��ڱ͊	만�~<q'l"U1��q@���[�.?���i�FW��2c�pv�GJ��X�iЈ����{@��m�-}�n���$����/�u�#I�(Q�ʮ���;)�ب[^2-CH6@�#J�|���)���l�����z��3(�iF�X,͓�Y�\���5ۗMbsg���H�8z	�\��3o�XW�S�O/r��R&J�*^!��d�0A��ź�Z��y��^H|��(��-�o��#�������Iᑽ� +���A�Sא�� ��~��Zws~��l'Aq:�����R��Ճ��)V�T�b&N֛����yce$�������Mx�
o7b§�.W~�6�:���r�Π%ښ9�����pi0JM�Q��z�6㱇~9,ٖG2��}�pܙ<=�u�4X���j�W��m���C��>��{�1(B�}�)��'M��/ٲ6��^�8LV��f �O��΋
�1lTǤT� :`���a���o������T7��V���jN�<��
z���o��T\�Qװ<��n �z
E��Ri��^�"�0�@��te<�Px�8�߸/��;`��l.}�dF�b�J⛮��3+�b]u��vGTs�ag�D�4Bs���<-F1h�=