XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ѳ����B�<Z�~5�����B[�bF+?
+1�[�Z�����©�9
&"�ߖ��,�N��E*�M�cf�$��� �N'E��n��]~u�ְ�cS�&���)���ϒ����ՂԧҮhIaߺO������Л�����a��YՅ٢���IJdm#�"��J�4��_z��Χ.��Ax0���Y���%-���)-;�D�1b��}gP�	s6D]�MF�~`��n�I�^C
��%T�i�n��*M�%����B�Ir��	ub������n��eh�o��Չ�t7�k�B�B��
(��c�6&ާ9<4���I�m|�|K�|�u+�<D̩��劃�������K/.����#�F�m^�^�:����T_�
B`��a���}H0��(�386�Tp�:Y1~�'f.�ɥ�'�vw�Kֽq�=�����e��U���1�րd��U׬?�H��>9E��8��R�"�|ߟ�������LuF����E~)zz�g�z�	�r@6��S���QL_KJ0�@��;F�Ѭ���k�"_��Nxzqʚ�IΜ�'{��Dc�s�}�K�G��c.��hK�D��;�2C�9�z��o+?�QY��ũ6���d�SZ�ك���a5ǩD
�0 �~�'|!s��1�+*��I��t3�a>� ��lk��u�43EJ�K�����yk�]0=ɻ��=��W�w��"Z�s��[������Ʋ����=��e	[�~��GO�J�x@�9%�\�;\�v]�F�zXlxVHYEB     400     190J��!�V��Tf�n/�k$sГ}u�Pҙ��,"^O��q>Pbs5��0vZ�LMo�gˈ��1�R	1RQ�;&u�/p�������(�]Xr �w�b�c�9%F_�-�n�J%a���f�����Ƶ_�ΐ�ح�e��u;)��ǥ�q�l).�\�,g\��Fp�/���wۖ��h�9���`�_��I��I�0�=�#"�*���ho�m�9�__�L*�����ƭ���$�8Ө��
5~������#�M>ӒB����2&�Y�yR5Ǧ�~�𜓦=�jF�Fi8�Gܫ�;�.����/��1�0�D�H�:�!ĵ܋���<f�w���j�]��G�*8�$*т\G�B<^W�>yJt@�JηM�IiĔ��6��~�=����`��_��R�uW�ζ�XlxVHYEB     400     180s�~Λ�.�	��2��i�ܢ�w�k�~_��y�`\��4L���5��U�� M5ߤ��(L�!�7�E�H�Ɉ��a�����
���8�u�:t�{IxIC�k�:��~��c��~]*����������$ːZ�=D�[J�Y�LG�5�n����C���e�M�{�5�Qvu�]0V=	�R��j�����X���4n�-�������m��R g9nd�v,U���b�pblġ�����2�����}�KH9Wj\���-C>Z%�ԏu�����g|�(��s��G�?�L՟��{�F�>�kS�r���	�8�lu�jb�ֽq$�LË�q�Y���NEMT��r�'��u�1�M
�nf�}`��rFϑ�dXlxVHYEB     400     190��������z��M��ܾ]�|o�\>5U��k���Q�=�"K`�@�6�J���NR�=���}tV>+����֗���%ո������*��G���$Jy�Β|οz�	�j �iMm����n_�gI��#��\r��B]|��	W���N����y�o�e(�����8;���ݲLБO�!�>�ʎ؃TC�+X�ځ,��
?m���5�s{�^-<{n�8�Mc�n(L��s�����&~P)��>>�q�Yq�w|� �HC�*��_k;��T!y�K�g�D[uF��@T���ʒΞ�.n�?�1ΞIII�8	B�;����M�'�96HT?�z�u�t����A�����)�nP:G���'��?T��05�[�g����try�:XlxVHYEB     400     170vr 
b�=g�w(׸�I��C4��Z�U;+m�:��2*5v�J&�.N4�zk���2�o�[t�����,�:�����/fe�m�6#���[�-���!��&��f�-��QC-�'=���m-�?�};b�l��<�a$�;�r��$�ڋc=ł��������#�_0ꥊN�F���DtY�`�f���VO�o������8V�#FLM�L�g�~�:^���%S�]��״�5|�F�s]_�(	��i���X�8�Y�lՓɯ
��.�X�!�vθ�5��ͽ�K;��̀j����ݞ"��X滋5��F���W�1�5�7�9�yt���D�L2{k�yA�q���W�w���~@��0����OJ������2�XlxVHYEB     400     1a0jJ]Ij�|A���.Z���}9����Ǜ���f[#��p���F�J?3�ƸKWdU����}і�,��h��׹�,�'��W]_��/5P>�S���n�y�����J\!��CS�W\8�l�Q��$7�e�[�x#�IQ�<ծ+\��D.�������I���6��7��ق��L9j.N����������c'�V�����@�LOf�IX<(��a��=��\et�-��u�:�$Z�,�AE*�QC����K�	��K[�M��A)���	����_�� jvK�e����a�!(O]�J�d
BHvp����
�w��
lä��40Qa/9F�W��e~���|�B�A��C�9��i��2�fH��yu1v Ί�i���c*.��s&���jA-:�#XsE$�E��XlxVHYEB     400     160$o�rܿ�HB^z���/�e�eL+ihK��� њ�3pu�-�JO�~�q��^�Yc�D�o�7Kځ��>�? �xYWЅ�e%O'��������O�30.�8<)�y"�a�3x�!�[&����xE|X3�,c]�<X7uڼ"�tǍ��Yd�ь��\�o]���Pș��_�O��Ms�#�Y���Ri��%�(�AJ^ڞCZU#i�svk+td����r��D`~�A;��˙��(~�$���Ѩ�V���2w)�z�]$5�z]��L�J�zd ���OT�X���K��=��W��JO�n��bnt�gL %ze}�A�;���7�y����%#�]�XlxVHYEB     400     130�O69N{h�e�����P[GQaO��Y�y[�,0�"���By�,�y�"b��ܰ��<U�A�@�_��<mf�������(/��#.�L�	��pΗ��ݖ�A��q���~��O�%9�67��9-?��a�?� %[rb�_�$V���]n�����r�0e�4�P�Xy ��2��j���Gs�ĺ�P����y�
"�4��I0����+/���PP]�szޢ��	���|���{C�')6�� 4O"�]6^a��X/�χ��>����_�B��t�Τ+	B?�C���? ��WSJ]XlxVHYEB     400     170|����O�F�h^���l��J�&oS
�. ��
���e$a���	����-��]���,��+�s~�ʀz!U�b��@2�n�5'r��V�Y� �ph�r����w�����yuKJ�F���K�]�!�՞�("s���Xr3p1&*a�v'�N�0� �,���&����C�#u.A�N���l�5&#L��cSJGcHY��MT��@�O*~�%���:��l���Q3���h��K{[5�q0�4��F�d�~��׋5�3�Z�V�������Fvn��|�a�J)��+��!�0Q�&���2!�.�ф�c��<�Y�=�v�ź0�W�(�����@W�_�z~1��$�ovk�܉PݷXlxVHYEB     400      d0�1DZ|h����4������*{�bU��Jg��RB�s����b��{��6Կ���g����(�\D@��*|D�
Xk!�2��It�N9��� �k����)�:�FN`�b@B�0^G.G6juY�i��Ag��N,���V��)�ʂ�N���k):[ǀe�aŦ�Dp���uo��+ϓBJc������j�Έ��=M�M=����XlxVHYEB     400     1a0��@Ue�Ɣ�'|Qاl�}�0' ������m�n^Ѿ��G��\�W	Ⅷ�R7Y\�<�t�X��Q|�V�Š���E�f(Q�R�	c	R�~�S����u
�]ք^E� �Y�����P�E,���^R��W��La�k�cx�z�&-`�+���i�^��|��9� 4ؙ�%9-�Lm�|�Ћ����aJ�{a���i�_���*�g)�]x� ɭ�n�>�)��L�s,�:�t2
{K�"v�� 	^�c:]�t\�K��B�X͞A#��Ao���ų]�G1,��f�u�I��d�-����|�U��%��RF����X}AM�h\z���\E�ڲp��O���ʞ��R�FnR����Q��9v�iMpCž`����$Ά��qp���G�m�ƭ�q��a��W��2
Έ�%XlxVHYEB     400     120�0lgr��sSh{�����J[����^��%Xփ��؀���e�n`ޯ�[�������Lp����pRژ��	�HJ/�����hP�I�T��b��P�49�a"�-�KH''|x����q�ń@e_0NR�1�K��ą�QO�Ԋ���� ����Rѱq{����p��@�<�ag�c��
 ��xB:L�bv��B�,Gv����~��w��$S��rݩ�%E�v�j�y���a�VSW
)�[�g�|��7�Hy�������`�MpX��
�ad�XlxVHYEB     400     170L��q��|�S=ු;r�F��SB�.��'�N���h����@�プ�-[� �Gm�w�]��vZ��%��>�J'��M9�gN"�D�F�4.v�����>����lCBa�)I��E�p5Ն����
}�[X�vY�?�ou�D���Y=?�;So����:��KJ�sA+?˺a;���k]�J<��/v�q�g�ŭ�m*0��3����v n�W5��XE�� fe�Fb�o��*���}-���f?��b��cB�FT��4����au����-�����'�VYy�2a�!!����w^I�Pm�����7����5<dU,��ի!���Š��}�zw�[(y��MJ������HKB�s�W�[7���[XlxVHYEB     400     170\z
0�.B"�l'�M�O��!���C�͛uQ��0,�fIޟ�A�܁�b�L���j�\g��EN��	�����9-Y��v��ޫ47�5���g�>�Ta<R����?�u�'�5�ў<��ͻ�E����������ӨA��Gr(�5\t��J�o����zX�=�����D��x��~�_N��֥h��w���¹@N�y�V��R�q	�͒��m��B���sW(1P��>H�Wso�����v#�̉*۬��%�*��N9 ����
�|������\'�R���Z�V	�I�#�~t#Tt��BH�������TP�y�*k.	^h��Cƃ�=��ik]����s[������!:���s?�BH��r�j�4XlxVHYEB     400     130��]@�QOa�sEb8�Aw�L�8*��i������mu�� �H�vC��,��,�+h�T���_D�؋���K�J1bpu�<�vR�/gVUHq�t�Oi֗��N-��	�M8���PAviL�[T,�	�ë́�3P@���,��q����8��W{�S`>5�����0���Rjm��J�U�Y�
t�����Y!܌�&�[�&�� ]�m�ϹMؠ���� 4���Ւ��ltN�U����_VYZ#���6	J�Ց���K���V��|Jj�7���B@^MY��f��q�phM�XlxVHYEB     400      c0��],����(�&=D��R�5�VE�>�[L�5Zusn^b��Ց�݁���s�`n��q��XƱ3�{�b��l�ЏtF-*Co�Ѯ�Gi�R��B ��2���mG�b9�ʩ
���D��1��E�uМ����ȕFE�R�7�2H���LD0�^u����j�}���߈4�V���)�>�$椐;�;XlxVHYEB     400     140'�钅�:�@��
�H
�&s��x8�Gʣ!�U��u:BQ��w!HN3xW�M�#��R��Wh0
�{���X~�=6N�����r�vBE��Z��0�0X9�j�g����O׊O~N�SX�!�vhʈD�D�H�����ةj��}���}�������=}����8t:�Y�������P�Ӈ��'�7��[*�+Lݎ�:�M�5!�g0�"n����J,/�ȝ��A4�jL���C
�5���1�U�~���DE�^��AaV�մ�b���GE�����m8���r�L~����8�L`����5�k�&pXlxVHYEB     400     160�T���>���F��LK�Lu��kb�����C�p�����ܢGVza&B�SyW�R���C���ϊ���i��z��6��ep?!+R]"�'I���#���R~�sZ�� ���|!�k�
ӷ�,���1�(HC~R�C>.΍��Q��+���hOa^n�!�>�`������,H~���F�]Z�a{7�B�� �� ����g���ɒ�G��>U���'Q�A�㐃�<K������l���Q����F��������;<�;��ȏ�x�ɸ6�`;���4��)H��	��� ��a�M��.5�Iĉ�3�`�e�%ɗ*�ףlC�E�]z��)�����=�GGXlxVHYEB     400     160�?���^�7�:6x��!�5�ZՐF�A!�z�e���ta���>ǔ��	����ivͺ�+X���ӕ�E����0G�
�E\�bqo~�cڒ�}�uۤ�]�U/�«�zϲ�g,A��Y4ύ ާC���#WXm���{�:v��5��:(@N����ܖ����\���ͅ܁�[o�;;��γף�L^����/��WNc���5Q�U��V9�o���I�M�q����S�� ��n�8jE�^4��-N�|�w�|4�t�@i3�����iϮ-��81��KOG!_�,\vWz�?'�x/V�c���A
1e�t#<���IeEZP�й�����׫�CТ�XlxVHYEB     400     160���2w�E}/��[��i�,[����w-�f�>���T��-�&���jJ0�Þ}d��e���TPZ!��(��ڀ��&�n��I�'K!�H싷����8tcE詓����wQ�7U���`	/L���H،ϙܑ_����k�W��8y��ѥo-��u"��zw;����Usk��Ю�]݇��1��n�Jto_�r�Y�v擘��rg"�=��D?d!/�j���Jk�Y��SPӧ�h[���ʆG6D��_b��4��� ɹo�w.����ßíJK3�(�}�w�Y]�f������,ʫ�VD0��a���İN_@_d��y���w���D��F���n���XlxVHYEB     400      80Ƹ��n"�C�|_l�٭�І&�,r�a%k�D�9Z/Br���	k� ��n�x%+�%��DmĝR��=~L&���ɴ%r�&M����9jK9��U�V\E��h~�H��	q�B}U�̒m�$2�U���XlxVHYEB     400     130�;(_t��� �t����܄��=�唼cu)�!8z��ơ�cXt�/X���9O�H���9$���҃��59�v�tjH[��+��]$ág�h�#�0&@�RbO�����Ʋ ��Bې^�����;\4_K�vu;!2�Z∔ɰ�DJ��΁�^�+�;��,�o�b�W�бM�r�/�h�.��2E5ƕ5X�@�?�Z��FV��(�V�k��&j��a���,�]�	���S2ݹ���v,5+߾��NI�Mç'dg���H�{Ľ�`�=�乓
+Ql4o�N%�b�u��XlxVHYEB     400     150x��`�/zg��0������Gq�jiÛΏ^)Ε�PJ/&K��5�,�ڹkD��5@e�?��
]�j��B.)mF��d6#
�@n��M���DF�VD�4��+^J{��\w|�$)�|!�}��K�2��@�@pL����5�������e�Ə*,E�^m��K���|f(��[<'>��>N�^@���^���Ȅ�銎=�+È�N�8�����d1�+��3�c]v� $��D5:��[�{?�Ǥ�q�0>c�����	�b�Q/{�@�q��D�.���>�.ڒ���T�)R�������g}��j�9�D�1*6��qF���(XlxVHYEB     400     100O�(]�ߓ�t&���T��ơN�҈��~A핵6��)/�.��h�튈��9�d�$&E�ax<V�z�O4.�d�ڱВ�2�A���!�zΊ�ſu��h4\9���@E�%�0RвpK5R|0�����
P�Qö�ũ� OJ}�6�&��<W������t7$� �s#�� ���U��`���1�AJ~�s �\g:>!�׀˼\X�n0��n�W�����^�[0҅��nWs<	���]� ��C����XlxVHYEB     400     120M�ã���3I�Q��d��}�ِ��ꂨ���~׀�g����˥�����I���@� ��'��8�pǽXoKl6x�c�f�P��g���Wɘ<6O��(I��~[?=�Jtl�0� �qY7��F�u@D��Y�A�u��F�2��`���f�$ݦğ� ��T��ʅL��_�"���P�i}#,��yk<��"�#m��5�p���FT؞(���q7�Ԉ�OaTz�l>��W'�(���pȚ:
k&Kz�Lo�~!�"���W��;��3M�s�� �u)�xXlxVHYEB     400     140gV���"w���P�Mc���)����iЎ�+�I����XB�B`.A/�a�-X�ute?�l���0�I߸���J��tx�U����c�R� ,����E&�e�@o8��C�嗣A=���ͩDu���=�!��l,2�`�+Z���`08�።_b6VY��O����DlS��W���v٩��.d�F�Ӭ?���@^q�XF}��/�7�ψ���b+/nl����û�4�P��~h�iQC/�����v�������ܿ@V�����, %�2���:�\'�sH}�Y�_���̤��-/�x9׎`.N��C��XlxVHYEB     400     130kq��6h�-Ϧ���U�aP�s�F< �� ��ʋZ!��j��є	���T�K����^	P����W}�����͸$t�h"niwj^g ����7�I�ߙM</���ao��\ �B��Əؿ��i�(�2gK�m6� '�8r���&�d�*FM��%�8?9�·�f؋Le;�F&�;'���W!֫�_P�Nx��e8k����J(O�"���|�W�^|<wy����a+D�[��g�?c�K�ʈ�.�`s'p�ʋ����(̹g��U����A`����pe_X�|�{�����XlxVHYEB     400     140���� �?ˈ6讀n(:�AQ>\��d,���ɠ���y9o�>lV+ߘ"�o�F�*�$�P�$A3l���y�߁8~--\�Pc/,�K��!cc���j��'vnI���:����2���Sog7���-r�祽���=�=�q=nVJ�]��1�AG����~GK��N�m�V���||w=H��޵�R: �=c�fV4�E1��9@%��3�(^8*�?��8�1z������҆s����l-�L�R�笂S�d&iDm����UM���U��H�2��2j֢a�ѕ�)���u�"DE�A)�o��. ��r���XlxVHYEB     400     120��Rle�n�Mv�&⬤ZE#i��v��?�q�&��Dٙl������(:�W����a�T4ɞ��.:͠�$!�s������ǿ�w {F<�㻵Y������e�\`3��I�f������K�K�l�L�a��R���ց�^7;Jw���h��8�؄h�.���3f��D̨�����ʑ%�$)�ֽ�פojud���6�z�7���sv���^����ZH�lJB�_nP=�y��K���9`x��͇�Ԅ%�bQ��^<b7��4I�o�X��DE�rJ�5XlxVHYEB     400     140W5!<n�H���7�&'�K����Z���g����h�j/x�#J����W{{Lc������ʉ�+ Z�Ц���r`�ӑ-N��?�3&�;+��E+H!�]�y�|숩e�h�f��B��j�67���R��QMfx� ��˯���Q�CE�@,�W�[���|��*X���M�jUjW�䚦ǧ �C���m�=k!J�朖��� �%4�s���NtJ��sՅوD�h������M�'����#��Z�,���3yb���񈳔����5"@�C�/>�ـ1��>8v]���+�~l� ep�C1�[;�Q�XlxVHYEB     400     140��P*c'"`�媝w���M{R����L��˽�tȨ��I	$�U@u�1B\`��#�ft :���Li�Qޕ3;t��A�b�]�)Y�[�g-J���]�DO�g��z%eX���+jx��GedW`�aw��a&�ץ�-i�|������1@m����3�-X~7��+P\�aP��{��ݖ��K�-~����ю�0�=v.Z�����fnRg��N���}_A�0��mx:����h�k�Jf��p�H�"G0�;n�ꇬ��75�������BcCG��l!b����I��>�\I�e7,�#5|k0��1XlxVHYEB     400     170����}��G���	λ
�L�v�k]��k�X�G�V0�����m�����j���]�}݈�MHǶ��Vh�����LX:�Ho�&�91Ckr�&�t�����{�m�R���xO�ð���Kw(M�Z���`8nN�
}����b��S��� ����)��vh5U�V���W�:�J�2�~�����G:�"�g�t,󬥩�z�(p���C|wV�|�d��k�c;����0��,ih���vr���t
�hwH�ʧ��;�;�ՠ#�]5㈁�t�P��	�0]�h��(��i�h�r���=���
�J鯸+,���h��N}MGKQ��Ȭ�	"�N��q>�m�{9�rM��f�T�qXlxVHYEB     400     100��M���K�?s�+�����ō2��EB�� ҟ̮pC?B�'4 �̀��9_{F���V��)3X*9�MV۶:$p'�ټ�|����}P�b�{�g�G������ck�"m�<}@ -���9���d�ۘ��c��=��������iÈ����G5~k�+��N4<v'h��T�So��5���-a��� í���$��W��D9Z",փ�%O���"J)p�^n�ƥ�r�p9�����p�fF�Q�XlxVHYEB     400     140 �Ul˵k���YTbCXB�|���������q|���zG�7HC%  A'����#&���튩�7�SG�wh�:���Sil$j`S�UkB�h;��۷�7����7�R�œ\���W?h@��Ep��N�X�8�ԍ����,���Bq�:!��M��i�g����#���Ъ �}�{
�_���.�~���B���J�c`����������
�0��-[�	���� BQ^�EcM!L�x�u˂�M�`�~"U-du��ڎڂd ]8(?VH��K�!5�7�ЄHZY�"�\��#��wvN�n~���UM`�!�6w#0�XlxVHYEB     400     130?J�0�)S�r�H��\������������Uk6�Zt�f�z��G�d���,�[�"i�^M4;�P̄����9��+"Ę��L�^�J4��������q#eAe�Ǔx�Ϯ)�j�S�y,#9����$���<H]�蔁��3�<[��^%8!u1ee)�a��3e�Lʎn�iԺ��Z�,��Ş�<v8B�kҶ��U^E��z{-������@��!2V)Y���?;49��_p�bq�:`��hB,"ܺ{���TZ歴�$����CR����#����4޹0��
��reD!I��*�XlxVHYEB     400     140���3�Q�6���߀�h[�+��XX{�MTF��9�ӳ��͛_2�t�x$���S�~-*�G1�Y�t�;h��4$�Pp�O/���g�1�}�"���.]/�Fz���V�4�H0�
��4g��Zh�6E���$��7(�2�!�)�$Ɣ��dZ��f��r$�@��`��>��_���K��x�wO82](��>;w��΁q���Cc=��+궫�9pzc���y��:�W�
.�|��xH�p`'S��!&Ä��?�];���3gX���VD�L�x����7�}�Q^Y�� F0>M�2XlxVHYEB      ac      60ߡ�/Y.� ~�K�E��A�US6��ȏ����$F��5��o)R\��*�k�)LϏ�����������F,������7���e��c!�T2=��Dl