XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190[�PQ{|�.2���߰�ÿ��G��
u���M�����x��k$9�����g96���v�!��{<����̫FÆ�HMھ1������&$��$�6m+;J�Y.�=���{=x�Ȝ��n�y\���p�7x��0P���x�8����i�(�[#��ҡ��_Ҕ'|�%�MN�����:���=O{�}gi�Xs�i�����"�G�XA����^��K���`�j�t~�Ζ��{*ic'L�5�A� o�jf6�92ǐ��{ᥒH>�W�"��=:�hM�3���p��E��Jn����~S�d?��G�������Ox�����Q���� WOb���,��L�D�1����L�d\�^(W��
ܨ	� mJQ��ip�s�|�G���ȝ˾XlxV61EB     400     130A��
'uؾk�Q^F�B�������8�&����K�C��ʚ�'�����1������E9�Y�#Z�������5����UI)>:���(8#�'�{[��)V��r�=�7�DOe+��h��y��m��#7zE=u�V��ݔ��O@������Xe�>�h��Gj�@=ϩ��y��&i��7��˴�D�dx��E���Y�N�S&�}��aV�o>�C�T4Ea�c�a8�u�nO��d�k�_/�؊%�IT�Z�n��[)��~��aȯ��N,Hj��W�ȸ,v�Ĥ�TO�,���=��$/u���)!���XlxV61EB     400     150$���Z[�b�l��e��b��x-!��̣R����Mf��ɐ���qƦ;��cQ�!���[�OX�i�xx:���z�0�t�5\i�D���`;���|���| ���73�[�8I�
.d�X��I��Q.l
�#d�d���x3kmr��e�����,��B���R�s��Hx/@��5R��^�"�kf��JS#�O,8�YOڎ����5�p��kT�|�x������{�Q�����X�U]�#MGpc}4c'v$��{�M���6��Tp(�$�Cdv��ە�%�/44J%��F�v��t��m����؉�r�_�"J��7?�XlxV61EB     400     140��_?�>��;�K�	�Dm���)��0C+�m���֦�. �����<N-�����.�ߔa���"����6�/���Eb��=�R���y�/�m+d�G��TK�_��Gg�+�ne���B���/�^�"����%?l�Je!nCD�"��;gX�b�G�l)�y�~��HJ�g��T���<��1},��
��l�"���O8��>��s*���)r=�g*���vޫ��O����^������Oҟ�"���W5�L?�K��!^S� �H�b0��᎜�'�LK^l�����V:�].��a��삎��t�k�2��iXlxV61EB     400     120�'ŀ}���(�'dn�{��5�Sy��".�Rm�{$d���B�Y�s�[_�b�&��g(��"�}|_���������}Ԅ���a� i��u_W|5aҎ��t=��[�.:>U�2Bq%���jw So�Hׂ:!�Z�U�+\0F%�ر�&�b�J�Nx�A�����8Rw��˰��Q���oB;�$e'r��*q��fݨ\�fC Y@Q�ޤ��,�\m�T�,��I]]�����/�\�$ǹ�:�v&ZR�X����"�ޅ�5��� lq��i$�XlxV61EB     400      f0��F'���F<86SQ���Ȥ�����z�;/���9kr:�kC�,�����4:T����@�/�	��&�\G&S�&\�1%A��I/ g6QS덨��۾+�|���-�Q�8}9R����6�-��X�����n}l�"����A̧�eٔc6�� ��ɐQ���KBk6s;
�/䟱��Ks�bk��O�E��k���s1�A�b\����K��R��Y:V�>���0�i��7XlxV61EB     400     120_���Ӈ0ߎRL�a�p�k��viw$�=�>�2��!�~���#k^}��g���
��^�2�%i����'������.H��@~�9�k)�S	�)"[�
���b::I�sX�a������.!f'��a���9���y,G �9�$X�F�<�	w�=�22w0#�J�f�F�!�ٻ!�[qt0:fc�VxhҘ4A���Z-� �%�MW�LP����Ik,S�w.χ_9M�����c��A2��d��F�9�=����tG��w��i�f��<B-�$�]��d�XlxV61EB     400     110���f����PG
2S��W�Fo�QI�y#�!�Kҧ����)�W|�	<�3�͋@X���� P+aƇ�(#Q�W�#n�a=��q�lU��ݎ���Y��x��e�$����W�y�ہV(X[^���(s�I7I�_肢�.��3��ٔM��	g�N�u����B�v�)�t>3�]�-�`�ԇ�0s�і4*y:��P�Q�N@�&�"Ȳ���?6���.%��v[�����d͵�mXҾ]����]1)e�k�����_ �y5��#����6BXlxV61EB     400      f0������̡=��qѰ�9�s��T���y5��耪�U�0æ�8��ؔ��cf���s�T>�oMo��y<l�0�52J���/�Xֆ��ЁeR��?��I�\�>-X�r��j�J�EougR�sz��J�w�>�҄)��k�8BіĽ���B����f9�	���~3�D���Mx��y�~��Q��7ǌo݂�v:-Y)���XU1S��D��K &�<�ʀ�a�,�%�@qKXlxV61EB     400     100%e�5��L�?/M����{K�.k�F�N�9���K��"��j�0��`�	]��K�sy��F8���pZp�3����R��^�\y�zߟ��B+0Fޟ�<��.���$�N8`|��>h�6��=�A�����+���N�nR��"��D�Y��b���i�L��m�Q����%��0�v��tj�2x����v$�~�r��8dp�:�Lb*�Kj�W���1���M6!I�j:�f�:��������P�XlxV61EB     400     170]�.���V�J���i��cq�x.���.۬�H�_�r[I¥	z�j�����=�9ΐ7�fn3��qd�Z�,��e����/&Ӑ�_v��2,�>2���a5�ډ]7r��u��������H:��� ��41�R	qL����2�]��
zl�oH������
坢Zа��]^�Yſ7�w�¿�& ��n������׵D[R���BL�:��7�K�Yv�ҸĴj� ��/{��g.7�?��z��³��2Qp�ju���5�-xb�Y+M�����%���@LEvzyu��Q8����Z��E����f]xZ����U_�-�!��%�Sa4R�7���Dj�Oi~�ժWn?�n�Ҽ��ˡ���XlxV61EB     400     140�T�9�!�+g���w*�TI�G�0��h�=���:��?�w�w��'��|�+�vl��3�
�ύ5X�͞xN0͚�(r����B�v�D�PM~Q� 
d���;��ר�l"D�N��
z�I�Ȓ \�Ԅ����Q3{f;��6vc0�o����F�.�MUp
Q�ߤ;I\��'{�ި��B�E������3ߧr*2���W��ET��j�p��؊��&�u�pK��k�:FZ�һ��J�g�:�;�K=3������l����9�z��Q�il�ά$��CI���z���͎��mpj�=ƨ��F��/p��X�o�XlxV61EB     400     130���*�x�����(����G,;�A{�8�6�nI#�ߢG��j���-}$�s/�E�g���s�&I5�w�%/����'��;�	SWa�f:RD��(ԁ`���۵��`����Y���'��͹�i��_�ֈ;JV�j?PHY�F��h�<��o%��>��5V�Wb��
�9 j��{u�깭� %��	��O�f|�Ĵ�'v�d^P;ک�_�?ݽ�i�4�?��r�z2�_���y�P��O=������܌���Xz:�Q�u�9�ejS��z�\LE��B�P�]#��*e��-���XlxV61EB     400     110*�>(W���p��#\yg���Te��+_n&�-4�r�g��$�F�α�s:�����H�,0pN��4�s.��y����_��Y��
�S��;6�j*����3��~�:H��A��Z���P�[���9��Br�o)���"�bU��E$����5y�tn��+'A�n�.W�ԣ��_)���Ъ�������������hz�*���Q[=�(�4��\���gV���0�l(�l��uHL@�R�b)g��.wrPϵn�$��%6��FXlxV61EB     400      f0����O%l��6h��Y����
�<~m�e��V��/�}ؚ>��g�$����.�lX0?IHx+��������i�&�Ͼ�#狔�j6Fj��k�ϖ5Zf�.f�e�)��i-M?Gfo-����gN���N�&ד���	�t�����`��|xE�jU����w�-�e?~�&ҙ�����ﴮ�u�L�s�gh�
!%�ioV����*�u>�K}ă�U_����XlxV61EB     400      c0�7�裈b��(�F�M� �����r��.� ���1�i	�p)u�^�d"���U�P��Bg��1Л�(�չe�į1	��Kw�V��$�W�n�M�������o7(���7[�`��*u�<�#2Ȟ�l�kՍ����;�Z���;"�Y�k���#k��'��ljL
��|1��Sj����<�1k�J�8XlxV61EB     400      d0J+���4m��D�v^�m�x���)��!�ü�WI:m�;��3���H.��i����8��B�A5d׆�#�:H�t�d��/�I���PKz��YIm�P���,��;'�������iۈO)ݒ��$��L�܄.%D_��}���U�~ X�l��'r��k��8ۣX�sX��v�*���S�&=�����2i!�)����5p�B1��kFXlxV61EB     400     100�C\�U7��^��� 货ѐ��������:�^0G~r��w2�噳@��f��GG[k�Z�1��-᠆s�ڙĊh���b5��%��ؤ���=�y|����?���Ub��(6 �&�P(�ʜ7"<���&O�S�v?g<)&w��F"I�c���"��*�j4Q���y��<�s$l�NՐ�e�SD��=/��r�O�AP�/��Ձ�%��U;ڵ�3���!�g�K�df�;C��K�v$�<�XlxV61EB     400     160���e���H����.B?�CK�v?"�LbhEǐ/MX��U��|��:&/�a��@�?�=;A#󿬆�́���͖��7�����H��4Bͨ�Kq%�U�{Ҳg6��oQ(�+�L_T��(�VAV�ȣ�Mb�����
Av�H�ĩ#g[�%�%D%as�o�B8@p��m*q�=!b+����:�����e�V���3��n�m��R*��}��A�=+���!h�v�9�`�����_��4� ������gWa%����ͫ�����7�:�A<��Ik\��mo��}��2�<8m���RM%]����ʴƳAT���PX������q��+Ȋ��ړm��M��DO�zw>�:�>XlxV61EB     400     1109�ZE�ڹw���E\_�cχ�O�����G����)Ꞧ�	d�x�R�/ѵm�iɠ�Q�Uzš�!��k� �1	24��8F�����f�P�����M-����>9.���[*����&������#�����G>�!`ƹL����0V�������8����w<�hؠ2gofT��U]�B��U�ʒ�2p
���Oz�����l�,�Bݭp �Y$���ǲ9D�^Ԋ�.����5g֥�YKN����@��+�N�XlxV61EB     400      f0�	5ԃ0�>�����x�K�d�أ 2v�?j
�Y��d�Ԏ�+k2���2�,�.�C��nyѡ��6|��h���V�:�%�c��3�OQ9Y	��� p������X������;�1�p>��"{��h�w�vi�A Y�^\[Oiίaݡ�qkgI*V�ygow���ͫ�\�J^�UORg@�vX�#L� ��
���4R8�޻g��(�l�k��<�H���e��PUG۵�	��
a��"���XlxV61EB     400     150"+P�6�W�C���%��2{� $(�X:�.�G��*����PW��c���%$�^�����2:>�=JK�B_f��O��h��dy�̡P=���^�r%�Iڲ|2���É�Po�|�����G�f��RQ};�d���́�u-�1��4��2D�2�.�5�(�5�6����ڢ�͸(�E!4w���e�W�u>����|�aDd�J�������������v�,>v����sB��t��>M����#�Y�];fA�u�:@q���E�a��0����ʋ@�X:E��?�X��	��ƻ��4�n�q?trLi�Q�(Bc3�Ș���;XlxV61EB     400     110�Rܗ&�l��{�Pe���Atۑ=��_��4澷x��@�]\2��^��o�0$; -"YZbP�ʙ��3q���Y}B�xU2	e��g)��Ͷ4J���t:Q�iá�����?t�+��&_�5<�4[��0��^��b�x׸���*I,�}T�ց�D]���,#���y>�4����j�<�h�&���:��2L<xI/"�'H$�H�K��
I��,�m���@Q��h%��"��.������o!�1K���?�+����H������d�XlxV61EB     400     110�ur1�[���~�C��Q%�/�y�@�5YEj\.'"ѣ���Ř�[,�;Ӟ�4�B
 ;ґh�J;ng���cvP�XMi��>AŜŕ�������sZD��on��Q�2��LW@������W�%9gU��(
@�$��#�Z��@�C�FHײ�o�Eo�t6Ӏ��H�s�xI�V<�BŘ>�c�S�����K�>ڃ''981�*�:#%�Ai&k"[>C���ǃ]L�ԝT�Bи����N�+&�a4�b�x�� F*V��TXlxV61EB     400     130w;�V�$*3I�G~��*~�
�\�u��+'U�dSM��n<����IeApa���ߢ=��5�?�ytN)�dE'-0���G�,�{�C�:HS�O�]�yam$EoJ�Ύg� K8��u"�
��Jr]Z�w^�c|@Q�꒖�b>����3�WV����.��* >�\1�$�n��&!��of��ts��QFd�+��7o���`m9�
�����<��]�9$5���PA	l)uwÄ�u����|�	�a���{��n�t͐D��[�^5���Y-5����Nk,��ɚ��!�o�h�GK��=�~OXlxV61EB     400     170���5���Y|t�9ֲ(���) P)�[{�ş�MR�݈�Wz)ϦD,���z�a��n'i`ej��0oj�<�q��i�6$gX�����d�?���X�Zu���rlk�L�Ţ����;�u|�y�����e+�Ci�
p�7���郄�C�d�F�b����vW�Y"���Wbɯ���!
�zFq�s���r��4HkR�e�)ƣ�\�����5A�UH�P||����@ RR������x��љ
l�M��oE~Χ�;&��n�T'"@���+9j�W:>Q ��K��1�Z�a�;_<]��J@Y�_oW�O�q�D���V^S`k�^R��L�k�x�;}��qF�2
��ҊH�*{�S�XlxV61EB     400     110	���&阎��q�k*JPv`>S�������u�K|��@���r���wBUL}�9�[gAa�)-R�?��UL����ᕡ:k �߈݃�� 8�w8��ݘ���\*NA_BU��I�����A<�2�2��tj�鸴u�NB�z-u�yen��n��ʩwؖmv��f��{�z�K"ia��}�S���+�.0�%���� A~����Z�@|*��������9
�A�r�XĬ���**u��?�$XlxV61EB     400     180��
`u"I
|���T��y� 	.3X|J�.�;����]P��шA���
��'���4f��Մ�m0���Ծ�WTڐD,�&rδ���+E\=]3��
@�ɦÍJ�K�C�M�£j.����^<�o v���׏^�eM�é����i�>S=nT���I0M}�Q�4�u�?�6>Նj������;!�����������r�U����xO	#էT�*2��p��.W�F �Oz25����k"���Ԑ�:"�vI��a*��U=�>R�q؄�_���m��
�+_���M�y�[�ff�T��Y��f��T���xA�=�Pi�Egd���@���#�+��5�����`����d I����ц� �jE��^�XlxV61EB     400      f0s�c�UG6|�a�q=��-5�35;Lm6�ey^��Y�9q�h�ȷ��F�8Q�'����AU2,/ytK��{�zh@�/2� d([�	��p{��mY2��u>&L����SM#\h�ij�u]�e����=.��9Qϊ�|0xjc�N�i?�kܤȏ�%�CP��^m����<0�t��*']UN�x���A��#��7_���$�
�=�����[��@�˰��>�ޒ�)
��R�k��XlxV61EB     400     110��r��]��B�aՃ�,�d���:��K�L7�V����m�PUd��$�cz��p�~�nm����l�"����Y�X�=�	6@����g��>:�1E���]��( ��T4rN۰bY��<�q����@���t�<>��e]M��t�Z/�A2���f��@Ծ;�va&���k�V�D�_�����W�ޠ���y��뎱�_�;cP6Bx�>*f	D�����<��t��|>�`)G�
R�sg�pÇ?,,��rߵ1��ƴ9�oC{(XlxV61EB     400     110�c	*y��e��y�ٽ?�z���k�n`qhDA��f3�d5#
�W��G�*��rx�u�lS-l��˚��%ĺQ�K'���EY�4��5e�Ф���p���-�a(���.:x�Ej�L:�y���qL�vc�R�&�]��hְ7�k���'��.'�%���#ы2�7,���c�tF'���L`j�hJY�����p�/ԉ�һfS|��Pʺ!#֊�=l�F#sC�lƁT9���d�s<~���۷xM�
��`�ѝ�~���XlxV61EB     400     180����lQ��$�\���K� M*f)�Ȟs�w��ʕ��-92���/���y�`��ڦ�Տ��Q�s3��.�՘�cPP�,^z�T��s�\	.��L�*�q�7���=�e�
LܲZ@�Y�U	��JJ��s���N�D�L��{� @c��(�c�09Wa��!~JV)�7�m�U��z������:r�;�/*�5��6�H+����j�8	 �e]�(�h�|���2����ȱ�O�~�/��7��*���M/S��E��ٻ���(A|�#�[b�����D����������`e[�Y���9>����W��c������*��1 K}K�DaHC0|� 2�*�{�9�d�f��-XlxV61EB     400     150��9�q����B�����&~���P���m2"�&�̇��������rq�f]�2�zef;�����$*���1�n�q��=b-w{UML�ݎv�W�v]h���!�~���QU�aΌ�?�� ��P���n����$�8�^}^�C>X�~���� ��m�d�d�I ��w�a�)�,C�\�����6��%E���76�zQ�F�B�r_��p#S�n����~C�G7<�J������`n|Q��T��*�Fĵ�tB$�'�9Y����U�~�����$A�!P���k�a�h%K��_����rox�mЊY���
b�Q@ҵK#XlxV61EB     400     130�Є�]~L�����&ҥ&HK��!��.XVUb�N�r4����1M�Ϋ��d���0b��r�j�?±�ux�p��7a܀�B#WJp�4�%�5�K�4�@�JB.[o]����ٸ�4�W@ ]<��J�{�z��1x��~ڶ���i�x(�X����۳\L(�r�n�����K�����֡D��I�K�&G��A�{���	c<.-��K9F��~�Qn��~�������N�z�1�zUtHT�Ed&����+��0D�a�z�YGoM��`=�@~�4�Ɔp6Tu�-,�u�h w��iU��XlxV61EB     400     140du�z�{-��s}�N��}L.�An$�*V_k˾�v�ڱ�t�� u0�L�F�O~cȢB#~�@/h?#_16)���rԮ�i0T�(��aUψ$��~�6�����ӿ|�
IfX+��wP�߲ܺ�u��X
�i�7�N�^�}��)*���U���O{.�m`�#Z������������;Yl���O_X��賃�C֑wg�S� %=��*�D�Ot�4���?���6�Ӗ	�����	!xF�_[ߊ��Mta�'���ή�&!-�u���p����D�(�FF��呩��F,s��Q�.�x�a��%��A�XlxV61EB     400     140�C6��`!���ɧ����橷.�j�҉�5�n=���3��<5у�a&��e}�&��Kh�ɋi���"��P""`����'��P� ���l��@9�	�J>=Ð$�O���[J��ӻ ���-PZg�}�o����<�Ph��.�w�o,������<�Y{�<�$����AK"�.+B,ls�(��s�xX�r�Z�M�i`�U�1j I_{^4=�����N��uc�hK'3��"/�������s<0�?����ѣ �Sg̈́�PV ��ne�2�[$͸��2u���T�U�9vX��CnG���K�������XlxV61EB     400      c0�����Z�T�D���v���=��'�4j9����dp��-]��J�:�!�]*S���o��JY�w5=�j�I5�"^���!�o���W�ly�J㪌�R9�'����Ddx��H�"@Zm��Q�	�����i���͐�y�鯈��5��/�:��p��MI=ߨ�n-�(���?#BΰǤ�i��%?����z;vZXlxV61EB     400      f0=��8n*�qWZ"IX�$zi1ZX�W�88嫪=
�p�s@�MW�'@h�{'�&\�N�x�I�%�T�
�Jkp��L/�j��4��5��V��ņ��d���8��rL>�gRẃ��Ἦ�1�.Z��$��"��G�=Ep�Q�|�Y�7���}������/���"\�@
XJ�,�������F�M��Z�f�Ѝ�8�k�	/�
Sq���:�TO���Dlg���߄���XlxV61EB     400      f0�+���	�3=��`+[�:u��>�~ԥ@N�5�q���3v	�˗�������	��FI���/ƳՏ<�9GGac`\J�2��aS4%����_�5X��m��%�Ġ4"�	O��w(�Yg)L�<
ڜ��j/d~"{O��?q��N���k.� �y�K,D~O� �j�LݢS��&��L��h��АE�>���/�:`"��5�W
�~~�4��ˇC'��k�*��j�6�B�������W��XlxV61EB     400     120�k\�OOD)4S�ةԨ\$�.�Z�����>U��[T�<��oS�P e��D5eǙ��{3�LX�"&��q>И�����-����7�`�%�A8�+��P�ʈ���.�G��	��b�����@1���W%�z�y��#�� �r3�|��b^sJ������T�2n� 3L,p�w��^�q� /�x䁍'���V����8�eU��(��Ti\$���M���"�օ�icre�V�5�d�|��};1E��{�?��%��CWt!�1����"�c�ș�ք�OwXlxV61EB     400      d0\lpҦȎ�u	C|�#�u�5�ۍ�3;����?T�że��؊o���Ro� :�v����z ��x�#��dx��9����4-rwNG��D�Q(^�F���@�~���q��S@x�E��(F��m�+@ga˯w��˧�Q�D�Zq�| �����4*�	����_��*RBo2q�k��p�E�`��'l.*)�"��t�5�|�XlxV61EB     400     110A"�6|x�$�]��,M4��J[pt6а9x~Zev���qT�v O�w��GU[�X;;�ɏ&�+r��08��K�j�e���l���I~^)�k�>Uk����;����[��oI�8X;����I]F<T;����7�xx`������G/E�$K#��E$'��xo�Ƒ���'�s����z0?�x=�� ?G�pV��<�J�r�*�6ø��rFיe 0_uAآ���'B�����@�"ӱ�cW���?��N�1k-�G��3���SXlxV61EB     400     120���PJ�)�H±�
��c,.׍�y�ʆ(#B;�K�0g!D�N.�"�ɸ�p�Ǵ�d��_����w���'c�O���'8V�"�T7)�xK��b�G5i����1���p�YZ��C�wTz��B��,M���|�]+�ˁ�pEZ��y�q���{|&�D��
��ې�Q^�h-�^�������FgV'��C?�b�1e��GB�95�"�x��C1�M�T���ω`k��lSkG/
`��{�Z��dh	b��j���]��/_�����c7p!`	`�`ҡhXlxV61EB     400     1c0���Y��V�X��ܦ�r�=7�vv�ǳX����&|�^�?���/gh���m7���PU�{�c��^rQ�#��'E$�<-�l�ϼO�a��[z��r��s��� u�Zl+�.?Y���ݚ���8
�v��\">׏�ɪn�
�C^L�Y<��,Ӹk�#����\/Ѕ�g�5^�DN�;��n3F?l_�4�{���L�|�Đ�{������n55�'�rz�U�a(*o�G(�"��W!��9��4��;�#>����;�L����nدvpB��A����t||�Q�Ǎ��v���S/���U��e���i�Ș�WÛ�Ԣ���S�Z��.Ѵ���PD��w����.�d�x���Y��:�J�<
��L�r~.�W�_����j��Sm��s�>�(�!�PL�A�_i�=�Q��q@�+NrV�~qP�/���.�`�uQ�:yXlxV61EB     400     190nF	���"s��*n`��*Dv��r�Slvck!9�h�`.k	��)!
��Ѐ�t��hg����"G:���i7�C�5���iîx[wp��"Qg%8jeg�EЄMڐp���r��cd��~�IhO	����j68&�%h�Q������+c�����|��7����u�����2��oj�i賌��|C�SJ��P��>x�`�?�oAё�i���X?��f�������> �`�äq_r�L�S����-�$�zpN5�,�l{h�r���p�!f�`/�9g��4������w<0�[dY���;,D���ǫ�1IH�LY$�a��ކ�Ha�q#��A�7�q2�K]�yl2���x�4jۑT�I��8��o�e3&	G-��XlxV61EB     400      d0���k��dQ������ *��N9�B��������u	"a�I�e/����Pn�JZ����J&9�;�E*b�@��5�3k��,amGt��M�Ԅ����mŬ]IPMٯ�O��E�kn�������^���?�W�4�u,�� �9Y3��c[�g��Ř�T���$*��
�)!N���ʑqeͨ�.��:�s=^S���XlxV61EB     400     140»�[�03�=~�ؑ�"�i�!qK*�^c2�^8���`W�γ������<ۻu��?[�	Cˁ87�[�/������%�~I��:u�(Utu�+�u}���DI29a�p�ۥ���Y��'��Jwf�vEh�5�$��g�E��
[O��l<���$�x2)qD��� ���Z�%Jhn�f4�*�l+Y�����(������v�s�uƨ���NHq�� gK��ܽ����D	��'�(�������$�����-�W���&5h�߾�����#'�7z�G��ˌ�D�F�R���JXlxV61EB     400     150a]��H/�r�iu�=��-�R~AI�oS��|��;��6�K�6��vE$m�y4K�.��z.���T�b>��ˤ��w�uios�t>*�N�\�E��(�獫�^ӂ�[f<�TP���TƑ�r��_@̮ߞ�a�k�2����U�QK�{��)H������s*�����G����2$�c�.)����� ��U_
"Ev�X�}F��E�B������8�3�0�1*�O6��G/;�R=e��\�]ǟ+��"�{�E��w\��F��v�\O����D)ͻ���h����iQY���
� ��ng���F�g������B�/T�>�Ay�QXlxV61EB     400     150������к㠘m	�G�P���ɂu����l�c]�n�1�e>;�t�x�� �@�2�=#�G����?��z�˩J�������\<f�$���s�U�>��&�Ul���4�R9E��g��(�<T�fv��?:����%��@Ys� cӫwcb<޳;9L�ns�C?�0QOqfa��*y���Mӗ,'v��J"}��**h�mw����?�W�E�-IP'l�N�N=IfA�A����|�!��JY�;����c/>�J����f��-��'f[����0�'��ƃES��Ss�=�P�u,̚3u��` ]�-W��#�	XlxV61EB     400     140����F�e�VGBwf|�M\�_��<��8�ky�P�+1߾Y@*�����r�T��˜���Ψ�k�Y�sSK� {����� mZ��B����6?��|/%�3����gлT�H�h;���D`9#�(��M���K���Pq,D�b1�d�/I4\�;yh������ӑ{i��9�õ$��V%}���V�x��� ����O�r��YZ}?q��C�s����h,�8U�&:�e%�uM�s���䡻�6�U\�p��j���S#UH��b���h̄6�@W5�;� ��k�����W%�P����1�����4��t��4�XlxV61EB     400     180c�Ή1:��á�b�W���{�y�$���������񳦖�y�y����Oug�Yb1F��%��xk�ݬ����O^�T>��?��ݿ?};��
 2�T��� s���n!��1�\Z;�ڣ�E�Vw|Rj4����Ӎ�7s4Vlt՜G�� �RV�_�G|;r���J/e/��\m��D��T� ���h�h����)̱� ��On��`cƺ�N�������������?*�J�}�$ȫ�������NEY�� �(eD���:�*��p.��E�U���������H�՝q�u{r�4�Gt)�&��Hd
�L1Ɩ��M���sq�E��΂v֘A&��2�����Z9�K�A�6����
�é��XlxV61EB     400     140�����TY�M�m�q�\�̯Aa;�d�����^�!-�_1ˁ�pK�2i��Ǒ/1*�u?/��ھR�.O��^��óq��"��L߆RFצ�{7��q��y�FUO���i��r>��+6Foo�������ĸv��?u�}pB5cN!'k+�~�*s-�u��5�\��o[H#]!F"k�0��ć\(H'��8���F! ��Fe�[dGu:�h%�j
��j
ʜ�tr�'T9gs����ΗJ���5����j�f������x���@�C� A#����L:]u��V���U��22���\T��&%�XlxV61EB     400     180?Y|ms�I�vy�9����xHm�,�h�
m|q�V04�a;9���i��z7<q�y��6X�.�107�:����G��"��{�싻{�?��NA�i`�.Z�<�m�a�MyN����ML�!�����ՐQ�|'$�G�n-�9I�pU��Y��.,w�t�w@�3�Sݮ#�˻KA�TD6���w���������ܸc�~�7;z��̲t0��q3�ѓ"k���1v�B�}�����D0�E��������l���m�6�.Ϋ�P!^>n)؜���錓�D����~)G1��rF?[��%��2w�_��b�M|oXN��^H�}�q/]�3��1���t��8������1�/^(����ڋXlxV61EB     400     150n���$a�d�hHnE�?�rG�8�v�߉Y.2WW6��/duP�1��4�{�}����]Nn�$tx(		(�w�+�m�E�F�+��>}5��CG|h0#V��D�
/�L�h�za��߆�L�J$�,Ӓ�D���R�ɞZ?�:wB��.��jGH�n�W�������-�
yޱ� "�o�q}|s��+K�.*aܿ���Q�!�<,���ko����I髺ҾC#t����{��Q���,� ?�ohġ�^˭��/�3�L�@�} �㺺He���V~�oV!�Pѿ\y����t ��o�GD�{-���ѕD�e���G!�Nָ�w�`G�3s�XlxV61EB     400     170ƇƠ�b/�`ʩ0*��`'�_�珻
�J�5�.���~�0<����1L����蒼�S*f'��PnpvJ��vg�h4de�Ď�}� ��k}^h�C$X����E�O2�ܷG�s��锍�}!����;v��,�Q���M�Z�ƿ�2�#�W�Q���#�\Yr ��B� J�����cg�sΗ��V��o?�'�(8�Ep�o��ގ%=|�轓DOk�)�R�e��C�o>6�I�A6[ �����2v���Hg�� ��,��:��4>��X@��e�'�Z*az��<&[s�;QHw��W�g���WA)`��G@Fx%�~�7�?�@�LH���Z;{��>�j�y��frXlxV61EB     400     190��!� #X:J�Bc/B\.�t]}��H�s��<��?��Z@T9[��� �T*��q��17��	�j	`��C��Dw��E\}����M�X��l�S�z�"o���t�����m+d���b }�s<��a1�GI����($Q8(�>��PV�#�%ߏ�1����z��K�O��Nɹ��=�poN���q��{�B*n�`G%lච��å��E6kP��1�Y�9;{���gm�uuX��CI!��<���P�~�t���9�}�v�ʫ�?N#�~� �C�Ӏ��٫�U퍡�s �I��`����ݞ�͕-�'y��
\.�bN�cMk�I<�ԑ�Ԇ�����xk��2�n>4�B�}x��/^�[vxn8:}.ќ����R�]��XlxV61EB     400     1b0��ɠ[�N�E-�WasFܴ�'l0Ǭ����%�ɸy�ގ����v�����㉦+�{�V���2{g���邱���EI������+
+`CD�祅Մ��^�i����Ө��1�g���w������*�U%y��޴�p��1���F����������B<2G㾸�k�2��NTt��* I�L�T0��&�s�I��)��I����AwTO x�ӹ��:ٚ'�ު�,��F�f�Y���\���;kLOLTip�zr�!�êg�s�������P��>��Fj���uk[c!�Z�`a�����]�~����t�7�7����d5�����f$�$�����n�^��6���1 dv���TWݲK���^e���֤�1�RA����ms��;|f�3:�b�����nz�P~6XlxV61EB     400     180�Ypc+C��5�3h�ʸ@������p��z=F�N�\ڭH��$�h��)��Ocƫ� �Z����y�Z�3S{X�[D썘2�F|�Y7:k>Z������w�NS�FX��x�drE�`�ea϶ң�����O��:�Dz��h˴tp�֍V��pѰ�_%�|I��X��ȧ�쿆l��ҍ���FEj�YZ�#Iv�)L�ӴiA�,���&�	�^(�aV�h���7i���m(˕���?��a�Jr��&k.Z	�@.���bp� s��>����{��qf�p�
.��=)'�4���r?;r)�s���"*�&������!��:v�˳�׾�N@�A��AR.�co}T�5���"~�2;����0�S�z�oXlxV61EB     400     1b0Lӂ���6�V�e��!��k�A)/R|�/R�
(4J��a;������@�5@z]�Q�(�i�K���/%�X�L�Ǭ�A�TNQ��x�����,��6y#����GҢ���f�f�����}E����r��Ҟ�|HZ��x�3M��4X%e���S�&2���^a�V��~6z�[���]T-e�1�c'����v�k��	��nFF+#�N��4��M�m+ej*Ʒ�C����H6�̒6����毼ɍ{�Sw��p@78=+EM;��?�	��12��GC����iZ�A��@Ev!=�s�d�=_���h8��j��}�<��4�]�"]�*~c;ۛ9|�q^�����2 �:&B3�_O���nt?�ZI����{���`��F�㒾Rt(�Ԃ:�lL(��P#�e��𖣺X��XlxV61EB     400     140�΂��ϑ�O�7L|{�<b����+g��4��D�n��΁���3m����в��H�Ga<-��z7�+��^@�m��]�\��z����.��η�|L��C!
C,��w`%�1�&K9�����uϻ?��n$�ǌޖ�Y�fR��iyL{ٻH�9��~��Zxj��~�N+%
>$ഇ�z�IɌן�t�Ð>%����Ԃ��:||3�`�9ٝ�\���r� ,J{A�?�R6�=˄���xgۍQ�$�*鉤�3����R�R��(x2�?2������6r�,�l?iT��R�R�b���O/���[qo^P��N-�'�֡�*KqXlxV61EB     400     1c0�MPD-O��8�V%�Y.a���RZo:�Y+�4SӳS^@��/pO�Jm�o�)E��g��]I�p�������r�G��e�5eCQ��t1�:c��4^��j0�,�Y1/Ϸ�G>ކ�/�G�L�*��g��6ـ;aٳ�,�Y�ȧ)
�B��x�P�����2��c�
Z�Ŀ#w�+����S]��$�3s���W���3��޼�=[]�J8�HL�[m�#X����h#`�}���i0����&�w��y�\��Պ�=�z�"f�*4g��Wc�ۚ���D��kJ�����531�{ �5~d�ؾa�˼��� ;LBse�������TݾCY�)�)�`ą]aN ��g������0��b�^�3��gF�*����}*�X$8KǍىee�n����ꐃ�u�ȣ�׏�>v#PJ�<nʿX�bvKj,'G��I��XlxV61EB     400     1e0`
T8
���5ό�,��:���ϓ��7�ͳ�����t2�`���cV7�xb�M3Y^]��Y��<i�.okơT��s	ưN�7�4rw]�z$��:i�*���	J��ied� Pt����|�;�:X�M��~:�,�� ��\��{B�2,Di�^k�J��\�1Z&pD�;�=͝�E�L�$AY��"��:�jI���3EZ�&��)��T�{�ؕ��-@B�rW&�#��wV�]rg���������;��K� �8�&�
e9]�1Ee�T__(�R�78̻���@h�ݒ* {?N��jrZsD�9I���U�goc��kf����R�໾�:�`�m`� z��G����������3�H�7�z����^������\)�u��U��29�1�
qO��.����CAs��aA�@A���U׸�?��פ�S�Ԡ:��0�lj�����a�1`�S�z�ܸ��=��e=_�zXlxV61EB     400     140��L�1�v��u�EGE�H}�d���ǩ��c�zϫ�|��\{� ��}���ku��N7,s�,�m���ț�P��=���O��H?S�h��HM��>Ǩ�jN�_8G�!�\�@�m-Y�OJTk
�r����G�5��,�$TP�!�佉���/؂��t�D|�u�a��LRi�c."�X�v���,ue�gڿ���I|i��s1��_�|,�l[	��-(��� B.TSǻ��$G��@,�j�-\��|����`�����x��B��=�AL���M�̟+O�&g�_����p�S�+RZxgY�a]@y4^������XlxV61EB     400     180���;?�u�XO��t�F��a�=�^�R��	�/������0bj`�[�F�?�VqcY�R�}��v����7K"���k ��A�T�t̠�شo@�{�ƁSM|���=Y3!������� ��10Tkn����i��}ތ�c�3�g'�K��t2I��'D55n�-4e�v[��٥�t�Ն!�H��5����h�7��-;����2\�Dռ���.:�1�`�=����lD*�l�[x�x��b'bp,fP}��W�8Z�[[EG�}�r�h�:�����+��$�8��V�x�ڱi����ݚ���oB���=����p�y�ȿB|����z�>8���<�z�s��Q"�R-�������4�t9f�Reb�12�C�r�F���XlxV61EB     400     1c0}}3��~ۯ9�=�D���Qr��^�V9��&ܧ�/F&=t��l�u���f��_t�͗��ߐ�7�ҿ��j�����ƱUP�5��K�y��m ͋ބ"�<S�X ������}x�d��O�c����OL��'���9��9!?o�<� >�9�F�NBN�(n�bF��%+�9Ro#o�|[I'��tN�0^�~;R���A
.?��I&�؏��CT����{�?�G�%枯)R3\q�ؕ�w`���}�j�N�e.��\���+>���B�0g��U����h��p���]q=�.���/�Y~y�u�<�9-�Z�j����(����!ao�ϫS��r��l�o���e#�Q1<��$�w�%�Y<䖃X7�N���z�NfG�
��uu� i&o���� ?��>#m��pl���d�_�גxt�.�(����N����o��ӌXlxV61EB     400     120�/�<u���]��M9 ��)�X�!o��u� \��R`��J8�����^��1�>%7�j�2���V��%�,d(>��n�Ͻ�GE�XtlI�pt!"��R���=u��CW�3�1e���,�4O�T*�6������G������$���V0�!�2�f����@���1�ۂ�qh���<���& ����뤆,���_SX`�'���x�ܤͼ1��H���v�[��[��\p��à.�P���O���8��l��,QT Mbg���A��s�`����<]ꘟeXlxV61EB     400     140��S���?���`�Z��xb�Ѿ���߇�LF�t�"T��G�p�ԥ	�uj�I�*Kxm`a�.�J+��-�l �SG�s��l��{��S�L��Q���]��wy���{�Cg�y�ɨ�_y���7�5���%���<��>�I%A�������~p���yΤ.[!��Hb��r��x#�����젅*�
��ZoΆ��S�����0
2;y���~δ"�4B���v�=[kd��~���4�*�;
P��n3ݿ'Q����%#��2\5�<���UngC;~H���p��T�TM �i癙�N6d_5�>ܺ�`XlxV61EB     400     160]1A(la�!��'��v��=�FԄ�{C&7�)taFʇ����J�v�,���u�-�&E���ye�Lw���QU9[tei[Q���ӹ�����yn�oA��g�9�'9��|�i�S��gw�2=�z������g��٬{�e�D�4K���xS����%�O�LF�(�Ds*�]Æv�E�s���矧{��t2�{�9��(������f�ڏ]'GV�3�`_�ޒ�s��Y���R�b����6����E_I�)z��˝|������p�%E���Ԍ����7�oox]DhQFX�A�6�����Y�+1hn+�
�6��LRbu���&�V%����=5u��E�C	ƍ���XlxV61EB     400     110������]��J�샍��H*�
꧛E!��?�ʼ
�#���o�K�1w*�!@��O⅏V��;����T�Y��z�a����_Ż������D����CC���D���s��>��*C�N��r���̾�G Q�nx�\W��.�5;�]��R� X3ECxNZ;e5�`:��/�/���1�>��Fliw[#�V�/�6����c'&Ram�z�����s�Gy5H^��NP5�"�p���yCB�l�Y��ˀ_GR��'��XlxV61EB     369     160������yv/o�ЦC�T9KC�@x�:�a�u4vM%���Or�]�@�佷u�Q'�Ѷl�r.��a����8���t�ȡ��@-0���f�����o;j��j�i���M��1�b�-�7A�������2*x[O���I�z]�M6�r�b"j�r��q��o����˦�'K��I�6�����݅�)�?h�
�m�7�HT�a���/�o�̅���_�p���GOA���LQ}��yO�F�Z�Y�9��W�Q�DI�/�]���dR�#�s\`���!+k��;.��.�+
L~�Q$A��q�]����J���JY&�i��%�Rc�����/���"E[��͎�"�E��B��j��