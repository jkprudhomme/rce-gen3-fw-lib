XlxV61EB     400     130���v�������b��3�%>t�*N��mc�rR�`oD�n��ߵh�����"󦉈��L���EE��ޭ3Ҋ�9��"���G�a�]�����a3'&����i�7
��Q�3���ޣoEjt��IC��Ǳ�U�}�~%)��ˏ��%P ��ٜz�2��8_(Ǡs8� ��9�oP����ku&N��^v�~�i�{�gQ4��}	�TmB�Ȣ�H~p�˿�S�����*���V������A�/D��	���u@���iӮB�[lC\B%�.��hf6�|�oi.�+���Iod�����@��+�XlxV61EB     400     120� .����[4J�qT���G��`{��p �ť����8���� .$�VX
~^�^-*2�����R�=��z���|�o]@�w.�A��&;�0��(c32��E�]�-id@���g�M	m��m5���c'�s�������O��9����S��*^��rw]�`e����VMo�����E���1�c�|��"��n��q�LIS6���*���o�� 2 N�{�(���ؾu.�����d�GW�BW�!�����76 �d�8ϔe�|Bw1o���h0zbȟ�!ʚXlxV61EB     400     170#��M8{�(��Q(�"A���u��pMƇ}�4�����[��ar�ZD��q�96�Mh�B�Г]O`1�X���A�� `�c�j�4����E%��)��5�^��:?�CS*���M�B.��@�F�6k-����.�5�ݠ!KJP�4��Vt@o漭�DP@�n$�������*Vi���k��,4���:��ƚ:"�d�0�Y�dz��Bm�t���6��ԇ� X��קo�^B��t�$�U��\)��#$A���L�g���߼�����ft�R\��'��	C�`�+po�H���i:ڱ�t�f��Ļw<c�lGf�eV��wY���ՙ����u��� �v��~�@��ᇑ���޿�<,� 4��|)��XlxV61EB     400     140�h��~K��9��rG	|�A�]*���cͿ@Ts`��4�m���&�����¦_>\E^UU)q�4��� M�@�LnL�t�dCxt�ڕ�ߨ�wǤ��
7-EW��H�C�$��U���f�*t��.`����|��Y�)�x��NT;�@Ϸg�V��'4*�H�6���3ȉp~�eͺ)|��@��Y��.��t �8o��<�}q�p�V3�A ԜÓ��4P+� tD����+N¹��=W���2F]�����2<�%�rO�m��dF#�#q�ȶZ�����)hBx�oѳt�&U�� ���< ��=s���Өx��XlxV61EB     400      60
ʙ�ګW������`�bX9O�r��d� ��,U�=�	No�q9��:K�{/����Ϫ���
��]�m�Ac�!�<Sl�U��]fxkk#|�{G�~&XlxV61EB     400      60�2i ��f�'b܇�v��,m��H�S�܄~#_�&DKa�Ӌ���i�:OIN{�VF��Ł��ǾC��8�=��a�%!�
 �l~sXlxV61EB     400      80���ó<b�"�P�'��5d�����&/d~�]�Gf
�H��1��m�ρ�sF)�ࠆ\��w,��!����AiT[������ŕ_�4I�c�d�Ia�eZ�6|u^�?]F����ÒXlxV61EB     400      90�T��?���c�ߛ��7�t���6P�f �J�����Y�\j���Ty�'�oK���cBvѿ�PN�(��(T�^m���*�(����;���VdK�2�2**��0�d6�J"��PN?�PJh�)���噢x�7m~y�3���^XlxV61EB     400      90슐���]퍒-�Õ�>�#���J�YBV^R��a�N��fN���)�����9{؆1I+^�fA~0zxH��^v���<���/�+���M��7�gc/��!� �`�ZcU���|�����r����x���[�������w�>O&��XlxV61EB     400      d0�u*���oprl��������}��u���q�;��[��ո�v2{�j�|�T�~�wY��g�㪢ugڝ��yz�N��
�6N8% ���XO�ˏ3�u�A��5M.f�MX�v59���\?<*|ק�bgVO60�v~�"z�p!t��Yq)L�1Xx��p��rCHl ���,ŝ�E�i=���'�e)����#z�� �Ij�˻_�Q��d6XlxV61EB     400      90;G��m!b
�sCb�ݐP3	��Xr�k�����=�w�JH�xP�]�!�i�zeN��Lɠ|���a�y�l�;���V*����I$�UNa��!q�۬(`x�G�7N$���U��,Gl�<�g�l�8��?H�tm�f�w� ��(zXlxV61EB     400      80�#Q�ҝ�^�T��MP1`����J��Z+�-�����LȖ��|��PE�G����s��CKa剖�309�p����S�s���F�3׍P���E���g'M�c�uM��J��cM�15�0H[�z�`�5XlxV61EB     400      60"���3�}D�)!��*<~�[f�Q�(h��UQ����ae\ct�N�Q�j���m7�^�W~���u�/o��	��)2���Q7�eV7*�Տ)�$��;HXlxV61EB     400      506�'�	n$U]k3fGb�K��g�N�Es�U`�ΖT�].X^���N�|P�T��jj:�4��"v����A�T=v������XlxV61EB     400     150�hX�W���!�����D����4=�"٥[��KT���g�$�$H]��Kxj�����Sd]�1d7̌d���F8� ����Z�7��� �"gͮԡ���Ϫ/���ܳ�wy$�}!8�ܴ�wۍ&f��O���]8�cɋo��	ա(am�}	��Â�d��ww���$�!�M.m�`Պ`4UR:!���z��Liw��숹vm�8#������c��������IoI�$/�&,nP:E�1Jjn! �-�ŕ��߬Q�Z�u������[H���ޢ���(�V��i��?s��z8�h����|n�k����2�d�zXlxV61EB     400     140�wd�w�rn����44y�)?D��j��,f����=��HD�?�����'ߦ�{}���~��K���� ���G^��=��H+��>���2�[ŋ)e	G�,��(�J�2���V�55�n�L�!���;4�L�OyF׫�dy��%I�\A� ��M/������d
�$�U��9dlԓ�>��X��=[�.��p��	�����V���'|m�o��Bk�r͋�2e�3U�י���e9������n��|f���}{���J���n�x��3�#7���p�ӯ�f\�M�ǋG�f�A!�P[�gg\���K]u?EXlxV61EB     400     190�\�W�l������c��ܞ�"�a)纺<ח��J�L7�;g�Pn���
�S�WF`EѾբ$��qY	�X2?܊���q1�;�H����Y��Q���t������y�����3u��2g?����s����G%��%�L�K�KiiZ�g3�u���:���S��Հ��(�
u�F.!�U�*��8���m�,KV�g�'vY���n-���5�ևr���J�N�)�0�8����b[���3*]%��~>����M����gO(�ǫ�_YvgDi8St��m:���੕8�	;�x����k�o��� v[a�n��#��/h��MP��� �'@�u����z�O�8���b����9�����0v��+$e�z������#�`XlxV61EB     400     1a0��d�=�W�xcD�MI�7r�'4�F�ꉗ\(�v���Ń�]����L+w�4�OL>�=\���bI����31
�	��Iz�Ѽl��)���K����D{�؈9�d�mw#��{���p=;Y�P�NvG6D|�ߘ�#���S����Bʻ�����2B�C����k�
`����Vb��G�<�[b��GPjdUa<�i�*�-ev����%�
L~I��pQW�x����p'z�G���q@H�\y[�Ċ�S�0�[��vSJ���y��ğt���t���~bIz~�.����y��^{#8Q7����#w0����%��P20����s� ac���X	�x����eFX��)U}��8I���T��4!ʀ�K��H1��
�(��"v��ȳ�@5�m��d�& 95��bXlxV61EB     400     120����]>��4�0��^��n.`_��abi��Z���Q�]�.;O`�<�n2�Y5�9M�.���✸�t�כ��K9~[�f1��I9Ӷ���w
�B)c+/����t��Gf�����ONW3"ʭ�%"H��N���	�D;������0����v���	���d3^Y\�c,a⿏��3�3����uA��=���.���?�Z�O5��v�A鎌�iF���c���f��;q<�)E	�鑈χ�>�+��̟fO���Ċ���J�_&
�r�η�XlxV61EB     400     130����O;p#��X#�>��C;��%>Z�	yrh�ۆ���ok[#o���DT� 
6�X?�]�hP֜��Ȭr0w�k-s���hN�by)�=�P�sQ��}�i�#�#wUso����˃\d�@�-��R$"�w� �$j�h�F�uu�"	�uTΑ����K3rg�'�z�aG�����|7�F��Μ�]�����K4a���ek�r�Dj�Zॣ��~2al�x\p��7��Ҁi*��{+�臨+�~EKR1�1P���I�9A#?��AR�lݶ?����
�S#qf>�_9�~]`�'�rR1�w���a�XlxV61EB     400     170z�B̴���:�X����9�w��т�[" Tt�^���Ѡ�@e	��Z/�� \�-C�W��� Lbo�
e���%>3�1�&��ZMP���]��f�z����ܧ���3�y��3 F�̆����B)��C��K�������< �Ǐi[�8�.�О�^�S�(�oe�����B9~��EJ|�7�D�;����14�0N]0B�,�3�t�=l�#Y�@4�hbZ�1� e��:�R��r�S촛�����P�TW6�&����շ����)D��Tnٔ�@R�E[Xu7���0:`���bny�P_1�����jQ"�з����C�5�4k�lB�h�ݷ��8|�n�/��	C�Qf����"��XlxV61EB     400     150fhƧi9,��[���dqz���m�BX��%�mAw���_�ќ K)�x8eJݵm�Ə9ts���A��g���>K��e��#�ʯ�e�"�=�o����*~H���eCc@2� QLZ��汬U���w)��ڊ�3di��)�
!c�S�B*9��X�[��  $U�@�zc�fŉ���ǳ-���AD���w���O4�YX��\�7fN����v=�$@���/�C�d���<��Ա�	���-�o�S�B`���+:��EQ^�iD�aEĂ;���TJד��Oȧ=a�
"�~�  8iQ>|z<-�>�'�σ�^�Z/�XlxV61EB     400     170���2>I1�5���K)�DK�󦩘&q�t��$-�0-F����y���3���>��"�w��0�o��f�(E��/���B��Bv���4ٍ��hC�!Z��6���e�1L�O�<w��(��)�{����s��G)[�a��=�0v��X5p�NoxR�x־�mʝ쩻÷mޏ��^�A:Y�� ����]ιh����;�T�o?���yc20J&�F#�o�=df);n�bV���W.��X��1��;D��-��|L�X9�`]������*��zR��7���rY��"�F���O���C}Y++U+��x�k���ن��JtY�\ ���h���3�1V�\.ը ���O��O0c!�XlxV61EB     3ff     170�΅Qى�g�T�|k�Ļ���y��j�p�Y5��Z�>���g�e	<�Bz��3�{�7~�Nϼ�ե���[W��%��\IK�o+��{!sea�=okRF��eX��\�/�8`��^��؜>��Σ��''��NQjX4I�#�|�.�ׅR�.�
�e��@;[q�ஓp)���ߩ��	����b�ȕe!7�\v��j�=��X&Gw���+&,�/�������\n�z���ya������Q�:�`��}#/D6�߭@I��<4u?��^Ύ2�4'u����#,��
���_L�����3�oZV>�hO�"��3�Ҫ/�1LP��л:�^O�eT�S�<���myc���{ʬ��7t�