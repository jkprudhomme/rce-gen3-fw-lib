XlxV61EB     400     130���v�������b��䥰-j�lM�K&UR���~-�܃�M�۫��F*�ɱD�@��>;�y��*n.^7�'�'��S5��"�����u�����FYJ2h��yE��;-G��.��+-=Fm���{���@��!E6w
{���G�y�=�A"s���"qҰP-��*s	����;�7���݅f�Ś�c���5=�çi�A�A�T���twaf_�W�ME6�K��2h�d�L�(���;Op�0�"���u��,. ��t
��W��uP�
�Յ���Q%��(W��@*�b�s�+BXlxV61EB     400     190騬����-���4�_y�3|H����/z$�u=0)�۵ҽ��!��]b����*��sz�� sw���Ӷ�6jZ���8�Ԣ$ْD2�̾{��d��ei�.��-|�˟+eFx��*~��Y���ܵR:YS��Nnft:X�	����ʹ{�Q���w�]�h*�}WV>��*��"���/P�@m+Yv۾E�?]G��
qY%ahߩ�{��M[㦈�?���;�a���1�t�.�"��pr+���Te�eTF~��(j<IϷ�3ۙ;�#�ڊs�aD��|1)b��x�b�a�����|�la��4�� gK�p�וi���ǱA��DHN�� �XZ�k74%a��~.�ͽZ�03G$�Ze�:�/��	�͌� sPG��Y���P��I2p��XlxV61EB     400     150KOe	8�x�s���N��XK�79�$���ĕ���'�jQk����F�Y��!�O�t#A�)�#�V!:��l�|��}ⵡR�.��6g�ự�?_�I��/$U�x�9�CN�8���տ�HRus|����}���_,���a��t�s���qAB0�p~�i�hȁ$�@���VԮ"���y�Q�K �iSz� ���O�G��Ep��^��0 xS�Fؽ�+$s�RGu,|sw�}կ��8�&�1nq\����
��r��UHω���j��`��em#�Ƿʴ]�����z%C��Ҫ[�����}��	��%ߦI,ԀCu�Ɋ^D~a���5W$XlxV61EB     400     18079D�փ`Z"'�B���$����B�u s�N�z�N��W�c�|gǃ����AX�1Sb�ډ޺�,��q�<���se	�;dW��� �
�tmL`e���q�k<~̼����[X:<� ܬ.@tȻ�Q}8
�r��#�m�=W�h�K�S�i#?z]�����V\�{�j����NMҌ�凖���V�FC�e.�?�o�q֘�aLǲ@�ڣ<��ߟ��>�^��61�.%~\�΢��sE�	?��D�R4e��]w_A*9Xs�0l.��������zC�[��iI�ʨ2wtkKɏ��E3��+�h��c�E�Ҷ(�z�~��܋)�F�:�8�)���H�"��[�V�c����[�BK�>xV�>'f�XlxV61EB     400     130��jPi�v�u���� n#dYN߿yn�z������w�"�.�����B*f=^�������ˇz����A��N�-����(Ķ�Q(��[g��i�z�U�%Q���	���1�S��!Դ0�)-����x� ���1��)v��u��i�k�[F+N玾��o���"���w}q) �*����x�N��4��㢁Kx�4W§��xU)�C�.~s�.9{�6��MN�g0�o��;���׿1t"ko'X;��#�0�N Ϯwڴ<�8v�ۋ���<����h�X�0��i"sځ�h6�X�7��R�ÎXlxV61EB     400     110��c)����g��*�6*v�OM#����Կ最#�9�Cf�_k�#�H���xw��[����=���'%�<A�t���zd>zڈ�����o�UkC�S��-q���)�<��R��Ě�#�ӘT�ga�gp�W��������c<4%c���fX��+
�A|ׅ�����<KD��.m!I;�#�7�'*b���%C:��/y�����eRy0��r}pBXM��q}��l�<�p��">�Y�G���2�*�"W�K����33��^��~v>�XlxV61EB     400     150h6�b�;#g7����:�� V�e+�Ӌ��2&m¥Mu��/��.r���)��x����v�e�GD�G/i`�Û�����}�W���n���{N}�&у�6�B�8s��!A<wyM�k��'�@�o�]֔����XTM���~����%D����9Iל�h3D{�h4�#���"m�s��&�Ā�^�<ƹ��Ub��3�a"�e�6����?Η����.��"���m�$�šj���m�v>6uo�֗���"�8Y��@�o��}	���7�X�HaYB?b@x�]>��Xy�ٿ����l�c_D������!3����ߏ��s�a�XlxV61EB     2eb     140��Ղ�I;��զ�?.����R�v���J�t�;$P9kڻ���-�c%J�m3�^��dVH5v(S&��>
z��}�ڸxˣb��� 2����;s���zH� ����M5~�R��jG�4���g�4}|�Z��:�^����@�lt�]���f�Y�'�>O찃������v�j%��K��t-�>�l���Ms8j�>�2�>O�%03#�.~��;�V@�_�U[a��!x'}��$P��D��� X�9�=x������L�Z� �0��k+�
c���t�̭x��l��[����n]q���