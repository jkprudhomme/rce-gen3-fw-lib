XlxV64EB    c2c9    1e80��	�~O��p S��TbG�J-!�1��M�5��[^��i�e	�p�%�:�^�Mg���lzM�߉�Z�HQ�1
B��J|��4�Í}1�!6�~ͼ�`��:�i������c���+�����H��K��֯J��|��B��;�V�v�UƏC�k�%��g��Nf9��۶��p�ng?�>9�����K~ApK�`B��v���lBQry85�i�����V�p��_����uCn?�T�l�z��K�G���s�*������鶈�����,q�rX�FZ�JA�k���	6B�6��EQ^i�쓹��5l�'%�Lt��p���s,ݲ��+zT��)�02��z����K�*�����%�����n.Y����s3��&�]��zM��=�J������x�D�{��7$#y����.�+��f�~�i��B�E��R`b�z�,�7�1Ee0괔����T��N��+�jH$Ģ�E[��t�&��+Jwa ��ӀXs/e�����7�SV�G ��$ަ���I1{��L�#�X\���j�;ol~��I��'R��(���3�bo!��ߛK�_�ݺ������hk��,�>Ջy�xl�"�|������G�J# �� j�������.���P��D��W���[�ת6���--�A��H�e}g�*f���W?{/.H��Vm�3����0�N�HzS>������ʉ� ϩϳ�۽2"J���6DF�$)�럸6����a�)�!̀����6�t,"Om���ޞ�E�luШq_6���mv�f��hR���8㽮;�.��@�:�&צ1��0ˡ����	6��Ԭ+��Oi�tb�j��6Ȱ�Z�%q��+�3���ΘFjs����7r��:��bā`v"�����)��?�����2�|�^��2%V��[CR�1��hǛ�{h�Kv�]����ݘEǯS����u�׶4�#�=�'`TF��7�����_{6�ƉRyBu~�)����*o����LE�bJY��=~�[��+�>��$HV�j�8���'S׺��/Ҝ��@���j�0�^��4���}���(d�̿�,e��rp�x�*�wcz�����5}:xΥ��GN�6M�]j��g��IX{\n���Gs����E�G����ω3.گԢ�.[{ӽ?�G�3�l�Q�-)#�o.�!TQ�W�
�,m�L�������\a�3^ �\t����X�rcYf�Ge���=3e �?�.�,��!YI4�U������es�6��@��01�i6�"�����l�.�+<N�3�r�0?�Vj�P����?�h^?V�7��h�3�)����a�m������[�s�j�ڡ(g���+V�1�M�}:JY�!��*�G�?^ۧ�}IS�h`~��tp�ey|��1��*�ʦgt*�٣����&�~�$�ś�j��8}��Me�[7&PD������G��n]jt1�����T
A����^�	���>~5�9�L�����j�q�?Ӌa��N��9׈d/>�������"̉��-��}�^�v�Id-���V�T��hY��2mWA����V'Ro��$ڱ������:W���� g��Q�a�m�9����t�|�M����G���.i=("�W��8�teV��(Lrg��|�)#q���R>5���v?�����0���XYז0 ��]��9*��'���G�1��й��V�~ir�(�e��D�j��!ȷA�!�BbIa�����GY��+H�"�RT��T�͌��G�ov����
`�׬�ҡa�҆<���B��B��j��%kO���(�٬O�>;K��6��Vi"X
��>�ߧ�,x�`��`���&c����������r�HB���'��z��Z]�l�ϒ�ꕠ9:�-[�^���I�-���^U(83۸� -��5Y��G��b�W�	[�P�G̐ۦe%�mB��
�>�~=��`��.�/�_�q?��2=�0}i:��J;y���A?��L�Q�����x��G�r�jTp��{�Œ�'{�a�ψ���+B�ё��_���
q�%�gi�k �c���D=���^�#��G�LT9p{�u�V���zHU=4+���
���}����k�����
^vf'����߱����ʻ�yt}�S�9��Y��y��e�Z�P#�%���Q��F]��Wa��_�cԫp�*P+���Ϥ�3�&{�>ԣ[�����Ш�2?�!�=(�,*m��s}~���~*
;���Jk$d��zӵ>��J=���+�	�TUe��� ǀ[��V�`�%��Ͼo#��,�V ~�p��^|��0���4�#��S��eÓ7x����w*�KFkuq�--�3E�5R��$v��13�0No>x!5��6^4z���K�~F[���|�˷d�z	[[�d��=WE�^ۚ	���=rxf����R�<�J ��ƻ
5o��Z��X���v_W�)��V���u��.�'3���^nۦ��x8���{�֯� ]l/Iu�a�`{zeI(E�������^c���@�i�[c�lU{3�5�`q��˅�ex�����z���3�1��V���Pס6(�ZS�����U��@5CǦj�;��-�"��F����������E�����@(�w�`���P�Qw|)}kw��|*��E���8MP/_��7�S����1�/Y�ۗd���� 7�#��X�
@�b�ǳ���g'�%`dW�o�xDQ�\��>�4���u<�r�-�
�I�-G�"oM̋"��;��Ck�*6S���l��(�-It7�+WKAՏu�9��'j\�p�jo���-�N���V�_`e��kd_��3�Q�"����ƊPQ�H�G���\TYܩ�ï�	Dq~���o~%��;����$��(�YV*߷x.�J�pWk��uPjR��I$V���=�a�A�/
��v�v������}D�+�a���f]�(��6a��!�i���'�o�߆mw��bW���:x�U�H]���[^4O`����V�/c�F�#��t�����s:�\�9�"�'?� �hr0Û��C�:q��`�pWs="Dx�3録��t�	����ji	�W�{��d�6E)o
���0I[����0���ڭ���L����H�͞�n�t��`
���J��/�%tgo��z��Ĳ{�3���k���={Ƅ̾����u�y����3�k�I��?"c�$����'���
#��U{_@�S��q�/{�M�<�Y�^�-���w�㡟=i�I�� ���gƁ�A�q��18-a���%�`FfK{l�S��@vu�GȢ#��}(�L�ξ�� �V���0��r��ۖ
?�~x |Q��j_�*�Vn���=���1=uȫb�2���qW�'ϴ)����w��P�a�3�[a_�F,�SPXu@nmq���8�3����/�Χ��"�NPp3�AG�Ok�C@�m�RN+�*�X��Z��JY49�v~ �P�5H��og�BRT6j��ƍO��*��_�1��	G/Nx�#����^0��kh��(#��� -b�q?�C+��ƍ/�	�N��ŗoV-"}���nU�j/�%qS��3�$�O��֠i:�W�C{�/C���̇i�'tt����.�����:d��Vh&���v������#����[�f=KZ=�P����+ �,}��r���L�:v�������5 ]Or��ӯfC��!����n��<����"��a"�%�S��?}2
�<� � =�}�P��uxW=5Xf~Z�&�7q�����Y�L��>mF޸��������r�^H��o��1?ݚ24y��\w�y�[�1��)����聮DS^à�?E���c�YYs���ZW8�S�J����7��
Lܔcaگ�2y����	��`w��ã���ٷ�λt�������K\ʙv���ko� �s�F�%u�ys�
C�Tu����7Q��@�-�'Z�����T]1��~(�EcԻ�#}�m[�Tn�� z4����=VI�+�Қ�u�������C�ٙ�]Kr�]Q���r��E~��x���z�����bؓ������?��l��
uu�ߙ���D��'�1��.��mS�.\m^D�� CUjh����n��9�Y��
�N_D|��M�35��m$�V�,i�'{�
.K]/��˹���<�2\�5�}-�H�jN"���a�Ey!�9����В޿6��
��H�@dD���|ں	`����Yt�q�ǣ�D�aA6	q u�0�-�sBj�d�/;�bEa�����A	��Kkf4+�I`	�P�;-AkD�5�+'R��5c@��븊�=c.�ZOr�sv������+)��7�vt�\ۅγ�$�]�m%2vT0�
��'��&����N��ё.�CW�2
ni��ܭ����8ə�u�1u�����Pf�J ��C���ȱ-��G���rH-�i����]��[юǣB��Ւ��fֽ�I��c=�4u�HX��Ȗ�J��@VS�ρP�? 9١�s����Y�?���n����SwH�[a��<J���]2��4S���w�6�G�+��[7j�L�«����7�ﬅ$��;f ӓ&w�u}���{k� խ�g݈.��țV�P�ђ
 6F��1�x��ןǲ��ᅬ��Ep���	;����a���X�R1@t��U'�_��/��G�>���ـШ4*��Y��O�(���HF���sS٫�u�PD�����M6a�&�������k�;j4�nz[��ڄ���>��-A�����m�w����G`�y 9{�xi�*���q�w�o�ZN3����/�6�OB0]����x��n�j���|o�2�*W�����H�a�{�a�J�hx��.@F�E*T�_{E\F_�_���L�@�I
�� A���InY�υ�S.���oM��<���P�liQ�����;���6_5=�v�wu�]0[��֊�{
�o�W �E	����QJ�8�2.�2�Q��|������;�*LO���]#TiX^A�D�k��z�v��#O�R��|���{9��K�W�s#�Nl��9��?ּW׊e@	�-zVZ���._�cDᝅ�����@鎈?� �J>0�KeÈy��q�u�Zɝ�.;�de�/� Y��~Q*��� ��1Cs͒/�\3DF���K��3�U7̿.%Fp�������m����D�$�Q�v�S{���5�K]��N�� �9�`�h�(؇��_�"$4�˗��bR�����'�l�j�ߐy.�Q���e���bqo�s�ldcZFg���_�4C�7"�Y�O��Y���2����c�o�U�5���7j?����A��|��1�h�{?(l�Z�V��7*���Ͽ�a������ B���d`�t�%�ȊS�+��g��q�^�x�+)p6��cq4w�h3��Pd.w�$�l�Z �	��+>�몃^�#�.ܰn�L�"{5{s��`���&�B��Izrcpk�Z?�'I���]){mD��mLY
߅���J^��kW/��f��$�u��	F�v���xRPnm�E�欫�U��N5���1=�6qq"��uV�MG�(���l��,*<��t5�r!��L����I������V3�\���W̓�M����#C�y�`�ݨ4�ӌ��#���>��Y?
\��G��~�հhl5���{|S���q�Z0ꭗ�nݼ�\�.h����z�(�M1w����Z?k�(H�J��a�!����_�s���J?AV��6�Ϛ@	�o7J��!�Ó����Q�F�3��<8|Բ�b+�U����P&|����~e�MF(�k��⎝WKM�s���\��D� TP�� =�e������܉:�Yn%�z�Z����i�NJt�H��~�f,��((�~v���@m��A
��y�x
a=���p�e��otV�s۟[C��S��"��߰���ea؅�1�5��3g��]�Y�e�.�I��o��R��Png.��y!�0b7��w�<�^�z�<��q�X��y�0�R���Pbp����p`,��^�ۼʺ����"(R�/�Q�OɁu��8����A��* ���Z�3;�,$Ȅ�u���S�l���E	g��G�+rWJ��b�4�;�Y��I˝MEϯ6���攫S��_���h(H��t5'|L��~3hnW�~��S��1N��5y�!��]�3e�̴lp�a��jt_2��6��ݹ`q��R�N��kja��4�Z�tc`�@M'ٵ���T��(p�7NRK���)bRwZ�n�AI���� ��Um8��3�H����T�1W���;�_���ߓ�Qr�(���PID�&+ʇ��?DjH�O{�Q낞;E[�dSv,�cߺ�%�fqGL6�('���C��k���S��q/��X8R�ר��:�����E��1���<~��7����U�N_H�(�;��y37��w�i�b���\����u���H��{u>K��Q�/_L����dq{�:����V��4�tC���m'd�dRR��^��]�蒌wa����
�g�	�f.zO7���VX~_NL�gJ��q�:/�Y ��$��p�!�}�^L檠;:�V,��ܮ�b�2ՙ�s^(��Ni43��]#����4�=Vzm۶6�����]�����! >�6"ي�R���tލ�X�nO�[g�>��ŕ���.$b/Aj$�6��\���4ZTW��j�cj�a�1�>[	�[�P��o��O�6(Ȅ�-G@X ��@����[m��*R�Ǧ��!! ʱ�d5>$���T!ȸ;����I��os��uI���Y�0A
������+@��Ż�>�TH�	����������[�W���m�y-	�V�3ٌ-�Щ��"y���)~s�Y�,k`�W�{1*��G�N.	ܴ��1��o;d=�Zm��)='.������@jGQCu�
�7�dj� ۆ����=/|H'"��4�H��V+�.&*/ׄ�ݛ�v��"�?��^>��0��"Ŝw3��Z�=�1ļ��EWr�������7������w@`k��A�r�&�]��D�1�3
��M}zSD�0��0�I���~�r�@����R/�A��������j���uX*1�׈!�pW�1:�����J���T��0:ч��qݿ*�Z[.+�4��"/�,oO2����r��#��<e6m0�H���N�"��՗h�,�vVR
�\����
��rSr&�#Z5"-;g�C喚�v��c9R��N����g�	�3���s�a0�K��$������Zv��3T3ؑ`�&걘��\��jzw��t����<�b���p��5F0	C���Q-}���!�qA�R�?�s��5�$�������UX��iN��� I��)%2����;Ƨ�H�A������?��HS�]�`.�\\l�}N��X����H�
m�=@R�5@"��Tg ZA�m��=(A#���s=�B'-��������{����s�����o��~�l��>L�(�d�=�.["݇�����.��Ԇy��tuA�H�!M�l��ɿE��.��#n0�6-��{�3������k�}~�(��P��s�k��������,T
Z�ϝ�k