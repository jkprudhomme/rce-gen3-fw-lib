XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160�����\>�Ɖί��M�Z�}m$S�Q��?��$�!�2��.������q�+�P�M� �����/؏V{���I�#����(��Gt/q�r`��� �@Լx?YH�e&DuC.����o��8�7^�ʢ����(����8��q4�6�Z�f����yq$��P-���o��J5�c+��^�N� �`��j�X򝼌�Ý�߬�P��`J��ߑgb2��l�zv�fH�V^~$p�ϖ3������=������jḎ5<�����=�9h�~�U�
Og���M����Yc���)}�C:|����]!,��;`��e� Re��a~��9q �XlxV61EB     400     100P�yj>�a{��i ��I�F$
&Z8)l=묹r���%�јe���svfk�}�iE;{�b��0��θ�8y	+�K�сFN�W	����/�ut.>�$�v�8*�$'���J;T ?3G�y*��(29a+��	�M�'e�C��6����Z\AK:����=ھ ��1oA�-�%;�������;sʕ��72���H��u�Q�ZkG0�6�dm�3�%n7�ݵ�t|�����[��(o�\~��r�<�n�h��XlxV61EB     400     120�Du��(�!N8-JbRG��O�qr�A)��~�q��;�B+DcG6�m�5/�2V�;��Nf(���rƘ���27:#!�㯔퍕5�# :���*�	�Ph-�`J�eS7pxl���W�i�*N��?.���i$����5m��H��T�\<(� =2'o��Vb���tg���F�˽9�+��O���DpN���[Z(C�1�ᐕI���̃�� Jk��bC���?�^6qtA������ˏ���d�J
Ue��2]7��{�� ���j�d�w!u����4�	�����XlxV61EB     400     150� .JI �2�Y�6߅�'��Yϙ�\0>�,�l{d��C���,dő��m�7�&%
yI��G�;2ڷ?����C&��j�:��)��$�yC�T՞�Yi ����{j�=Qn�@?�K�����*ƾ�!�������![xxQ |/y̱��ϋ� :M@~�ك�|�0��H���p�V�Ė�=����I�x��|��17�I���%��u�8�r��sbAo<�8F�<�"E:)PX��]�gw�<GA2*,BJ�v�0a�G��w��ko���=��(K��B i|����C"�n��1�&}]��|���[����[��ά�G�M�F��ءYR�XlxV61EB     400     170:#��F��D���#�B2(x�U�Q���G�~b�k��9m�o��շhZ����`..�� �����!�u�>������d,�;��b�+�I�ɬ��jH�����$�[�y����;��� ��zނ�,�oܖy03jD���ܷ��Sw=����`�a��FM�V� �%S�����%�ӊ�����ٟ`
�bz@oԷ�E����ԲOx�9�vM5����S?`D�������x�Ck��Fm'I�̺Z�Zϯ�[�jΒ���ܫ�ɏ˭�p��bd^�|Q���'?����vz+���Uq�n�]����7]5�P#� ���pY��rW]�jH��	'�\	�؁k��x��XlxV61EB     400     120{:3^ L`�u�{������gM��b���w�T�0���ߺI�!���zεT���hI��.C�~��<E礤"����N��U�p�$��2����A�M���͸�Y-�U��_yB`��N�o�{Ҷ�𽓘��6L
[В���r����:E����HϛtS�C*#��S��%�Gn���V�G��=v��{W���sIR߷��x���t^��0���R�}��zi*/0��L��d~�N�:|d-�,��Ҿ�1�G�d��Ə,@4Pt�$�loøj�4�=�XlxV61EB     400     110K|ю���x�8Vأ���XH��e�*o���qj�18.R0k���r���/�����-0L����,vB��x���[f���԰����$���L$ES]�X�/��<�/GY� ch?F�? �c���CڥL]��F����Gi\k�<^�M�_�3J���RxK��y	��S\s�ơ�c/���]��fu�20?��R�ET6')��4X�a6�Z}E�x@N���m����zF�
N��a��ѝ��o�=c�؅'.*Nv_�L	��XlxV61EB     400      f0�
�9��w� ڥ�].y�ך�vs�H��I�f��f����_�.qa3�3R���߇�6@��@T	�*(nc���mU���GQ�&�wl�d-/YB�Đx/wao�8uu���m�~��ڃ��͵=n
_��1�%�A�)���{0s����0av�>
���i�JB,l�
� �E��i����N-�����5C�+�/	Ty5kR(��!�УA�slp0`�>��@���6�[g@�ۃ�
kχXlxV61EB     400      c0@�JM��{
Djt5�nB+U����5������g?8̗��b�.�A�S�~g�τ�c��z�����1">������R��)L���,�l}Э{p���v
�b+/[�KE �O^h�C8g�Y�42²`������WB�A���C�u����-���&M͖�viZ�UMq��7���n �f�y~�XlxV61EB     400      d0i��jV�nڇ$~����Ѕ}��	n?����ZG
�!���Ǫ
����`����(��}Wip�|����#{n'-]�7���f5*�`6B��˟��J���ƒ��f�3F�N=:٘�M1ɘO��yj��)�c�m��4l���9c�E����F�s��lU�5L���̑�wX���ș�N�#�j�23���A�RK���zD�|XlxV61EB     400     180x� �@�Հ{����JU߸��VAJo
�Ԋ�[a��J��k��@=�8(���{;�9"0�U����k�V�҃	`���uC����T�5`��Қ�g��O$�w��!�CM�E�pvw�y"Ψ�AF�w�hg.^7A4k��g�'�P�^4�/
������T����>W�T�;dXuRX�L+klwz�
VdS��w�[e+,�r/�#��5��}d�y�!��'K�E�f[��q5������1�&�?HOΪUۅW�1![��m��O��UaoA6���V���t��v�����6��<�K�3Ӛ� �Q5��Ɔ)/x�tx��n�y9q�}��}�&�w�V��[�߫:���#�Pԭ���C 7 "q�XlxV61EB     400     180ܓ�GDwZ����z�w�zb+x���7fL:��V	�Orƣ�l�T��܍�g�����Nݳ����Y�v��������t�2VqmR�8�``�mQ�/ɩ�z�kR�Y`�"*9KA�����Է�Y.�Ƽj�ǫs��}򣞿�ށ��2Q��D��<v~]�D(<�0'	A`Q�u����vkԣ��<�̈́��m*ُ��yK��@�dYo��SL�&@ �(�$ն��:�T�kQ���0������ٽA��-g�=�L@��&��l=Tw��M���[N��0A-Lw-��Q_dq1I��n�GtZ�^?pߦi�I�����Ȋ�]}!�GR���xI*��v��)97���$�\�0e*��gJ�@~��N�`YI��0��8^XlxV61EB     400     150Vb�=�*�_.����h��C�$!~О������37	
�ր�,��|�e��a������x.�[��1�6�*��D'=��K�	zzE� ��+��=_/]�8'BZ`�g�ghIg�8�1��c��M���~?ڂCo��9}���B>�G��c4q�;/ۧ�+��W�+�f��bYG��X��@�qh��k���Ua�oO��g�#��'��Yf�Y�A�,]�s7��(�5�e5��8Yf�7��жH��A�r�̮cr#>��x<C�Sx$ب��6 �o�حBn���
��Z�305\�!~�M���!j����lJ���ގ ���Q��3����1�۲a�XlxV61EB     400     170#����Z���#��Q6��HA>3&��kk��,]��y��K�sH��OȭΫ�U.�2���Z�i��Aљ�nV����T!����?��>�[��(CmnK˸��T��t!�_�<��L�	N}S<���]*T��k�ƠK4s?���n�Q��>nA�j'b����#���������r�ӎ5���E����ݖ��C��о�����{n
���8�l�.u���z�k�߻�Zd����D��v�\�u!�rR!�$��8��w|��D*���ms���g������}�7ۆڔ�0��֔�u�CB���w�ly /*2���袴iD�]}�:��U8q�cDAZ�b^{�t({�\���g��^�����XlxV61EB     400     1a0�X)r#������,+��J;�l�I �8�I�ʩ��m��;�g:���P��=�zLC����L޲����_ ��������?e�������x����a������8J�cT0h�(��#t�����Ο�8C7��+9�.tJ�������h��so��@RSh���.ʫcǓ�筂�քXn�w�S�o�� j�n�'⁣U�;��!6j�K��a*EtP�gSi��Űת(���j���\�#1}�@XMH� �߲�o�J	��EJ��k����tMVA��9������5}y�LG��o�[�,������N�ޕ�Z�:`��C�w��x#�z�Y2d:t1!ht@N#�՞�i�j�����T���|���dsW3`a�gRL�SM�8����	��V_N:�H�XlxV61EB     400      e0����FB_|*�t�C���iZ ��iے�>�v�^ν��¨��%'��Ѻ�U��VzM���&EJ�E��yܷBCZNM��L�7��4�@����%�H*3q�?���f���DuP�����ZcR��"��:ҺD��_P`�hB2C�ܨ�м�կ�#�M�>bOʓ&7���4`Iz8����.h╠��!�.��V)��0'K=���#b_�~g0�g�T�w��Ѡ�TXlxV61EB     400      f05�A�dR�n�X���E�|*o���-o�Yk��M�18-P�B��@�P;s�Ee:?�fJ! �)Me󹼝08m���A�=���vV�#$?Q@�Ε����}7k��B�|�n�̰��Az��
��T˖3�]�>�Q�;���il�q55�Xb����q� �ޟ'j|�,T�2ͬ.���0���"��ɸ/�ԟ&�Wx����f���䋊F3�誝�^D�r�3�p���eč5XlxV61EB     400     100XϚ�#��_�����d� ��Q���Erx��p^r�o��m��	@ڙ���^	r��""W�/#3�Y$�N��Ē5PE36�M�`�kލ{s���ҍs��G�H�B����*;�[{�G�U��J%.t�c@��)��t�Y��)��� ;����~4l�V����Z�h����*S��~���j�joL��\�
����:%��� �'�4ձ�]�J��<�.�\2Q����9�}�i�&��İ?�	�hBXlxV61EB     400      f0��#P��9�l�5q9D�!b�%��D�B�J���EMLx���\����J��u�$��uX����#��䚎�����E�=�%Z"�${�ኩ��R�xa\?��8��E����d�n��0\�_uǹ@�~�f��$���Y���܃��t��?H��)c��Z��<��'&N���{!��T=@]rcE�C ����t�J�L����ڙ\e�� �|���z�ݵ��?q �k�܁&Z�*��=��.��XlxV61EB     400      f0���;��b�~Բ��Ja;߰���XI 壴��� �D��O���k[�.�p��w��/�v���M�~�~�uy}.;�����s4/ Ԛ�L]��!��G�����_�L��M
65Ǧ�d��r�Z��y���)X����Z�3j��&Po�%K��(b2�h���D:V9N5�ㄯ�����;�el{�ռt�}�&�5W�F�<���)��F# W�/7vU�n�#6ia G'XlxV61EB     400     100f#�,�G���٩��/!��$��q� �z:��S[�ʆ,@���H_��I&�\��;B�mlSoFP%h��J����|r��P�6�*�o��@}��XVlz�j�a��8@�S�����?���`�>�e�Rďx�%��������{��8����'2ӷ�i�a3��?e���#�?l8��Aj@]F]%I��l�ׂ�w���K���^'�oM�'!�߇4/pۛ�O�%�#���AB�O^]����e�"ɅXlxV61EB      a1      70�'�U���g@�Wk�*�����|Pf�Hrǚ�i���:@㩱�\xY�E(�%g�oCT��b����������mHx*��|F�[��mU�޹d��B6� ���X���eU��