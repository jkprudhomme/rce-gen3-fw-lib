XlxV61EB     400     130���v�������b��䥰-j�lM�K&UR���~-�܃�M�۫��F*�ɱD�@��>;�y��*n.^7�'�'��S5��"�����u�����FYJ2h��yE��;-G��.��+-=Fm���{���@��!E6w
{���G�y�=�A"s���"qҰP-��*s	����;�7���݅f�Ś�c���5=�çi�A�A�T���twaf_�W�ME6�K��2h�d�L�(���;Op�0�"���u��,. ��t
��W��uP�
�Յ���Q%��(W��@*�b�s�+BXlxV61EB     400     170�_>@�a�e�z�O{���f�$����q6%Mָa�|�a��G���+�ע�K����g���/f������#�&ȣ��Y�N`�f��F_�n��#�LQe+׏�sQ��3I�v�f�jd��$-���]o|VDu�	$�;��J4~�|��<&����	�W(����~���rC�;����@=8���zK�P�<��h����g"����d�����e�,Ƅ2���.�T}�u���.U9"��F��z;E��b��5�ϕ�:{m�j��=�.h"�Í�U�ƀ�f�W���W-;?��E><�{�$�P7BV{ԆDC��2��[�$�Hv�w�� u�A���	M�)بa��j�[Zt��,�0{�XlxV61EB     400      f0�4a�����K�Ж֢
��A�ax�;�#BR�6�@��[�hɐ����rʫΖM�Q���9 �W�?B2N��Ι
F�ޗ���̋M��3�H���6VA���(�� �t��Vah:~�ＥM�qC�W�"x'9���_/���=@�N
����5
����Ua��u>�^�$^-��,��ż��K[r��j3ZgYpY!˽]�(X��T	k1|�׸R�\�*tR0XlxV61EB     400     140	��J��5��MW(��Wc`�k�P��d�u�u~��7-�i�����#�{��Atx����
⓯)VUv��	�;>�4vj�s"���	��#�X'��-���a͸�¾��`%f���6po3��\�b�V���i��w4����
 �y��+.���H�/�Eu�X>�Zf?KT:�ZaBB�Rpa�=c�.u�	�%ڋ]W8��t���J���
<qT� �H��n�~/^%��֑3���V�(o�]��3�y������V4\��EtnJ#�����Q��A����*f����+�</e�"��i���@��#�ݽ�XlxV61EB     400     190�*'5l�s����{!N)9ŝ�6$���>�Q&����	���%�UO7�/`M����%e�LC{�J�GT�K���
+'��&���F�?cg~����I���iG�@\����]{E
��l��뗮^!İt��r��H�
^|$k�!���j�f����.��t�^>ހ�.%8�3��R9?������+�dVI�3v�ET(%��Ic�0]}����?��C���Ӛ�%��B�+O�9�vrT��l{R��#+T��,��O�n�g��:`U�5R��2����-�;���H��*��f����sxY�T��L\����vi����&tf:4��k��;����A&�#z��/H��̗�cvZ��"��[o�%�l��_Ȅ��{�'�����e��ߕ��"+��XlxV61EB     400     190_(�-�8��Myޚ>%��Ui�⟹���#0���.����XQ}�)#A��6%�����|a������a��!���'�e�3��zuQr2��tY>��'JN����Yx�~��6�uFOV1�z�V��Z|��LsY>ÙM�6��
��qMU�W�ҦɈ�����2Cq@ϓ��:|ّ2锛�̿�� g�}>�T���T�
��ϴLR���@�T����Rk��~�0(_�L��ǈ*dC+t7G���a:l�l ������0����Ò��@�H��^�>jЊ�ć���J��o@/
0�O~�f�Gd-�ZG}��(�*n|.���jG�O+�5��,�w�.U/ڃt����D�d8E��fޠ���2�jȆ�Ъ���ܛ�����ҝ�id4�ඳ*89x
83�}XlxV61EB     400      f0�U�Ь7�ӹ,�Zc���
*э!����ɩ^�|¥"+� �%��z��x��qg�P��H��Z�-��8CU�K�%����J"
��;'�sE&D^qv�e�FS5��Ǡ%g�q �cu<d0��m�ɷ�;L�sJY�i�4���{��3#e�w��ꬎK�i��R7�*^��;�3>��,[8&3GÝ%E��!Gw��8���Q곏����r0��hÖ�8���XlxV61EB     400     130^���x��,��|i�W`����G��#����_���h�QE�\����u�)\��t$n$XY��q��?�JA'�E\�#�\E��8ڦ��L�Q��$��[�%oqk�2����`{���4r��%q����Dh��߱3s��?����㧫
+8��_���#3_h�V�?�G	t�������t׳�i��b�R�K<�אѩ����Iv-E�m�ي*��ރЊ��A��j*P�p�X]��Pe:t�$tB��9"h)��XI�zu�hL���W�XK� �9J���P{���6k9�E�XlxV61EB     400     100��%*�ʹ�r�	8ᱥ�EUu�2bA���1�r���o���J�@���Q��>���؋���C>���Sʾ�_L؞��A��>�%~Pma�$o!�bb�JQ~���
r��UӔ�~Nͫ��<A
F��q!�J���`���ҫ"�wد�=�X���3&X���I9"���� %גO�hv��WR�G�j�����x<�c�\y�?���V�� ������X�Gp���C��[�`�����A��XlxV61EB     400     120zi�l`�	�aK�u6N�����d��SĀ�K��G�Q�0W�[":�9�ə��w���k����da���Ĳ�ۉ޳��������f=L�ꃎ�{�<������b��Q"Se�<�����06�;�2��Na��I�!��!��xv{����	��!>�	�W���G�:��[G�����	��Br6�� ���~��-x���,=�����q��ƒ
�R�[�&T��'�N5�+������.���Λd��B�>	�Q���i;U�h$��o%��Z>���jxXlxV61EB     201      90��!X�97\0�5��p|�;3�������d���p�1�RgC�|XH>;�-}�"��l�{���_��P�*@��8��[f�6�٧�@t�B�MѦ�&~2,~����C�����}9�z���䈰��.wi�