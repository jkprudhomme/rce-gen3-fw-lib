XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a04Ll�k�Ci����i���0��+��s������Ot=a7�'���>o��Վ��³*&�oi�$&H�L�jZ3Bg�z7WЦ(]'<�w,�Ԕ~*n�7Y��%���B��z���rǐ$�+��M�L�0�	�Ri5l�=�)�s��/X��Ä��u�.��8��; ��G��@[� ���^��r�t#��s$��%��?��Y���:al��`�ā��E&�ňl��ǈ�t{Yr� վ�m� ����|J`����[�"Ԧ��pl�-��/-@qp�i3
���2��>�O	�T���?�jIS{�{a1ڨ���W��ϥh�I@���T�͙��Ks����+������S�獝P�,�s8B�&nQV[~\X".��:v�����ӃGXlxV61EB     400     180���8P���U!��Lf�$�p�ڭD�#�U�-���5bBî:��m��na��>�	���7�R!zyy�X=��ۺ�^���*�W�b�uG�"�37v�����FFHƒ6'��;:џgÂ�f����r�V�m�Oc��yI�Jt�'j:B��]I-�� �}=��F�[_��iB�Czi�$�3	r(�K�pg�'V�:�K��a+;D�O�ypݏbj��g��ظ>m�0�+���'؊Ĳ��UI?��R�B9���S"a�G\�Ăk�P`��8M�`qq�\��nÊ�8~^��Rk� M�|r�a@#k�i=g3�*��2_��q�֥��ݛEI0��H8K箊�ެ���q��9�O6S�jןP>C2W�(KIXlxV61EB     400     110O=�UT��a��D@Z��찫��f)n�ȫ�lBX:v�]XFo������u�_��g���)�=y�Q�ƀ�g�r�{H�kGw��S ����_����-�0z�EX�m��7�k���tjc�.�+X{�� �oj"�k�;s�䦱d��H���__yV�eO@g:�a��w'�9�{E7C�a�l'��_��_
hM���`v��9t��$ϒ���`�� <��5]ֺ��&M5��b�����	#���a��1�ʨ÷�XlxV61EB     400     170,�d�b!Q\�0`a���a�;� ��s���4��H���/�Ɛ�H�,}��b���~C����qj��Y�q93-]{C�\�VB'�y�K�MzpA���5�S�W�ܜNB{�OS=M1�M�Ϻ揞9@ŔL#��l��ao"Q�0��0�x��A"�Ul
�ī������- ���!9�u0�"?f��p���>����v&.S?�
�q���`�llc�_#�V<:3�Ew-�,���!���gI����:.��s��@<Pu�29ٴ����,w��g]�<b�$9� 2�?g_U��Knr���=ҕ��I�|����F	:�T�_leBi�3k9�Ҥ�ŭք���[tG�z���%hϖw��OC.$�8.,XlxV61EB     400     140yM��&G��/�'���qT���������"��&7���߳���	�]ڌ����7�����Q��H�@�?���|���2c3�	�z4�'�[p����l!��:kB��㰶!^�Q�S#�<}��Bl��lѿ����ț�_�I�n ��`E���;�C��tw E"��V�EC���f�O��flęT��z]���	64�.��P�s�Ɖj�%f����IE	���>ԝׅ�;>j�����!%�4w��鞂t$�S)�ֿ�W��V�J�ʹU��#��%��)�s��\W�kH,~���'E�[͒f��>��. I��XlxV61EB     400     170��*4Ӣ�w�z���S�\�[A�I�o��cR��NC�s��9r��c6��� �\���������"O}�آ[��@����>����rs'.FY�~��Bl��Sd��yl�X�yX��/h�?�Y��ba(q�P���Ȳ�v!�O�Nr��i #�r(��[k�m�?��1��%��e�j1?�9��]�4���-�8��7�U:��=D�Is�%��yK��S�I]'Pv�oHĨYz���HƓH
�.<�g�q�|���%���������{'������F���W9lH�q@����u������RyL�?�d��Kܜi�W#4C0�6� K��|�s���ZY�Kh����>������qn^�NXlxV61EB     400     150���>s}a!�vЌ�d^���'�Y5<��� a\�p�W{+���_OZ=,�#�[�i��V�=j���LK��(�b�ӆ9���Õ�9.�'!��{Y�����v%j��-��f�c&�#�1)�!`K��s�M~D������T�.��q���lEj�;Y��!�o�~��a�#��?��Lڳ�i *S��jln���s�����ɓ�i����uү��~8� �Y�Ƃ��8��09a�� ��o<ej�2�qW�|���!��]~jB$~��ᒜwu���k ?�n�(�,�6�gVCa,{���%��TK�(�4'����x�0�T14na�HU�db�?�.XlxV61EB     400     180��9'�� q1�r�����i'1@�8��J������`�#��=�����ɠ?�M(~�c�I�������|����2� ZE�h���c>H���#%P�R��D2�24��q���R�eD���A��)����/�8Q���]E:nx�iɊ��!w�<����|��*��7��a��ʚ��4$4$���B��3���^˹��N�Y�~$���=��y]'n-������a �M3�ǉ�UE�6Xp*�N��H�k��J)���t7[6q0Q��u��_���~ņCjPs�j���8O*�_!� ��F�f��q2g.�uMjO�rd]w���T�5���(��b�߉x)�:�H��0;�4rC3u|~��5�.�XlxV61EB     400     170tl �eВE�y. ���|����OB���\k��<ӝ�|}+��5.M���) J�c������Z��E���������U,1��C6��P\�oa�8�ʛ�b����R�4�Y��7�b{�5
�O:��A��o�Y�w`0��Ue�<��*Q������g��!N�^n뿥���a�?�2��0��,g�`r� ��T���gKg%�U��Nl����HR�w$n�G��QSB$~��D������=�z$gr�Cȟ�W���������9v�'Q:}�M�
�U 
T1���7P��!��+lH�L��B/�,0����b��?��S�Ϗ��}<�}�ˬ�Fg��nMa)�핿!�^:(�,d1�-XlxV61EB     400     140�@�{n���S ��8Q��h�Ae�������{�F\1�k�icWyR��_5���=���W��q/}��������
c9�wh��G��P��/A�+i�ͪ� ��MNv}�.���gB�g��W����� C_����X(������Yg���`;!�}� �)��gW�W68�����C�vy|(�e�+*PᑇW�4q�p��8�⌤a
�����8JG���ܛ��q@�|���!����c��5Y�5Ѫ���<�rDu]�jD~��Ƹ0R$T����ˎ?M��d��2���<�j3�-&�C����D�LFXlxV61EB     400     140��&R)��K㔲J�d�����"�&�af0��.dԯ�ڜ4I��G,������>sN"R������@����u���v?l^"�oE�7�Uo����0���I�!f�2m���u��y���,����j�5�,ѕ��Ja�E&����MEJ`_7�}��n���J�.�x��u��Ut\�'�j�u}�XJ���Z�I�,���;WDZu��})S���AYy2��%+EEB��拆ڤ�����1	MiE� s�&r2.|���Ե����(��U ��b].Q���3�|�Ÿ�Z�q��%T'&tu̘~����jD�&o�XlxV61EB     3d0     120wK�Y����N�IF���w��(<6Kfpg�a.��a���k�-�޸�����	院4Æ:uGh�=�I�9��wL'���K �#F��g�#�N �YGp�(s���+��(��QG��8���ΪzYv@��G�Ow؊�9^�k{��K�y0��LGd+��gLѦ�3�f�M�-~�i@!�Tk�LW�B������{�Y4�6:pP��q��hr��w�����+d��,Ն��re{���~�-�Qv��zf�mG
\ȹ�a��O|O�JO�U�C��3��Z��Q