-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.2
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : zynq_xaui_gt_wrapper.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module zynq_xaui_gt_wrapper (a GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity zynq_xaui_gt_wrapper is
generic
(
    QPLL_FBDIV_TOP                 : integer  := 40;

    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     := "false";        -- Set to "true" to speed up sim reset
    RX_DFE_KL_CFG2_IN               : bit_vector :=  X"3010D90C";
    PMA_RSV_IN                      : bit_vector :=  x"00018480";
    SIM_VERSION                     : string     := "4.0"

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y12)
    --____________________________CHANNEL PORTS________________________________
    ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    GT0_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    GT0_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT0_TXPD_IN                             : in   std_logic_vector(1 downto 0);    
    ------------------------------- Receive Ports ------------------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GT0_RXCHANBONDSEQ_OUT                   : out  std_logic;
    GT0_RXCHBONDEN_IN                       : in   std_logic;
    GT0_RXCHBONDI_IN                        : in   std_logic_vector(4 downto 0);
    GT0_RXCHBONDLEVEL_IN                    : in   std_logic_vector(2 downto 0);
    GT0_RXCHBONDMASTER_IN                   : in   std_logic;
    GT0_RXCHBONDO_OUT                       : out  std_logic_vector(4 downto 0);
    GT0_RXCHBONDSLAVE_IN                    : in   std_logic;
    ------------------- Receive Ports - Channel Bonding Ports  -----------------
    GT0_RXCHANISALIGNED_OUT                 : out  std_logic;
    GT0_RXCHANREALIGN_OUT                   : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GT0_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GT0_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT0_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT0_RXCOMMADET_OUT                      : out  std_logic;
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GT0_RXPRBSCNTRESET_IN                   : in   std_logic;
    GT0_RXPRBSERR_OUT                       : out  std_logic;
    GT0_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - RX Data Path interface -----------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT0_RXOUTCLK_OUT                        : out  std_logic;    
    GT0_RXPCSRESET_IN                       : in   std_logic;
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GT0_GTXRXN_IN                           : in   std_logic;
    GT0_GTXRXP_IN                           : in   std_logic;
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    GT0_RXELECIDLE_OUT                      : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GT0_RXBUFRESET_IN                       : in   std_logic;
    GT0_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    GT0_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
    GT0_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);    
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT0_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    GT0_TXDLYEN_IN                          : in   std_logic;
    GT0_TXDLYSRESET_IN                      : in   std_logic;
    GT0_TXDLYSRESETDONE_OUT                 : out  std_logic;
    GT0_TXPHALIGN_IN                        : in   std_logic;
    GT0_TXPHALIGNDONE_OUT                   : out  std_logic;
    GT0_TXPHALIGNEN_IN                      : in   std_logic;
    GT0_TXPHDLYRESET_IN                     : in   std_logic;
    GT0_TXPHINIT_IN                         : in   std_logic;
    GT0_TXPHINITDONE_OUT                    : out  std_logic;    
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT0_TXPCSRESET_IN                       : in   std_logic;
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTXTXN_OUT                          : out  std_logic;
    GT0_GTXTXP_OUT                          : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GT0_TXRESETDONE_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GT0_TXPRBSFORCEERR_IN                   : in   std_logic;
    GT0_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GT0_TXELECIDLE_IN                       : in   std_logic;

    --GT1  (X0Y13)
    --____________________________CHANNEL PORTS________________________________
    ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT1_DRPCLK_IN                           : in   std_logic;
    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT1_DRPEN_IN                            : in   std_logic;
    GT1_DRPRDY_OUT                          : out  std_logic;
    GT1_DRPWE_IN                            : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    GT1_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    GT1_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT1_TXPD_IN                             : in   std_logic_vector(1 downto 0);        
    ------------------------------- Receive Ports ------------------------------
    GT1_RXUSERRDY_IN                        : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GT1_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT1_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GT1_RXCHANBONDSEQ_OUT                   : out  std_logic;
    GT1_RXCHBONDEN_IN                       : in   std_logic;
    GT1_RXCHBONDI_IN                        : in   std_logic_vector(4 downto 0);
    GT1_RXCHBONDLEVEL_IN                    : in   std_logic_vector(2 downto 0);
    GT1_RXCHBONDMASTER_IN                   : in   std_logic;
    GT1_RXCHBONDO_OUT                       : out  std_logic_vector(4 downto 0);
    GT1_RXCHBONDSLAVE_IN                    : in   std_logic;
    ------------------- Receive Ports - Channel Bonding Ports  -----------------
    GT1_RXCHANISALIGNED_OUT                 : out  std_logic;
    GT1_RXCHANREALIGN_OUT                   : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GT1_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GT1_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT1_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT1_RXCOMMADET_OUT                      : out  std_logic;
    GT1_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT1_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GT1_RXPRBSCNTRESET_IN                   : in   std_logic;
    GT1_RXPRBSERR_OUT                       : out  std_logic;
    GT1_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - RX Data Path interface -----------------
    GT1_GTRXRESET_IN                        : in   std_logic;
    GT1_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT1_RXOUTCLK_OUT                        : out  std_logic;    
    GT1_RXPCSRESET_IN                       : in   std_logic;
    GT1_RXUSRCLK_IN                         : in   std_logic;
    GT1_RXUSRCLK2_IN                        : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GT1_GTXRXN_IN                           : in   std_logic;
    GT1_GTXRXP_IN                           : in   std_logic;
    GT1_RXCDRLOCK_OUT                       : out  std_logic;
    GT1_RXELECIDLE_OUT                      : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GT1_RXBUFRESET_IN                       : in   std_logic;
    GT1_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GT1_RXRESETDONE_OUT                     : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    GT1_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
    GT1_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);    
    GT1_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT1_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    GT1_TXDLYEN_IN                          : in   std_logic;
    GT1_TXDLYSRESET_IN                      : in   std_logic;
    GT1_TXDLYSRESETDONE_OUT                 : out  std_logic;
    GT1_TXPHALIGN_IN                        : in   std_logic;
    GT1_TXPHALIGNDONE_OUT                   : out  std_logic;
    GT1_TXPHALIGNEN_IN                      : in   std_logic;
    GT1_TXPHDLYRESET_IN                     : in   std_logic;
    GT1_TXPHINIT_IN                         : in   std_logic;
    GT1_TXPHINITDONE_OUT                    : out  std_logic;    
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT1_GTTXRESET_IN                        : in   std_logic;
    GT1_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    GT1_TXOUTCLK_OUT                        : out  std_logic;
    GT1_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT1_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT1_TXPCSRESET_IN                       : in   std_logic;
    GT1_TXUSRCLK_IN                         : in   std_logic;
    GT1_TXUSRCLK2_IN                        : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT1_GTXTXN_OUT                          : out  std_logic;
    GT1_GTXTXP_OUT                          : out  std_logic;    
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GT1_TXRESETDONE_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GT1_TXPRBSFORCEERR_IN                   : in   std_logic;
    GT1_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GT1_TXELECIDLE_IN                       : in   std_logic;

    --GT2  (X0Y14)
    --____________________________CHANNEL PORTS________________________________
    ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT2_DRPCLK_IN                           : in   std_logic;
    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT2_DRPEN_IN                            : in   std_logic;
    GT2_DRPRDY_OUT                          : out  std_logic;
    GT2_DRPWE_IN                            : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    GT2_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    GT2_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT2_TXPD_IN                             : in   std_logic_vector(1 downto 0);        
    ------------------------------- Receive Ports ------------------------------
    GT2_RXUSERRDY_IN                        : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GT2_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT2_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GT2_RXCHANBONDSEQ_OUT                   : out  std_logic;
    GT2_RXCHBONDEN_IN                       : in   std_logic;
    GT2_RXCHBONDI_IN                        : in   std_logic_vector(4 downto 0);
    GT2_RXCHBONDLEVEL_IN                    : in   std_logic_vector(2 downto 0);
    GT2_RXCHBONDMASTER_IN                   : in   std_logic;
    GT2_RXCHBONDO_OUT                       : out  std_logic_vector(4 downto 0);
    GT2_RXCHBONDSLAVE_IN                    : in   std_logic;
    ------------------- Receive Ports - Channel Bonding Ports  -----------------
    GT2_RXCHANISALIGNED_OUT                 : out  std_logic;
    GT2_RXCHANREALIGN_OUT                   : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GT2_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GT2_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT2_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT2_RXCOMMADET_OUT                      : out  std_logic;
    GT2_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT2_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GT2_RXPRBSCNTRESET_IN                   : in   std_logic;
    GT2_RXPRBSERR_OUT                       : out  std_logic;
    GT2_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - RX Data Path interface -----------------
    GT2_GTRXRESET_IN                        : in   std_logic;
    GT2_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT2_RXOUTCLK_OUT                        : out  std_logic;    
    GT2_RXPCSRESET_IN                       : in   std_logic;
    GT2_RXUSRCLK_IN                         : in   std_logic;
    GT2_RXUSRCLK2_IN                        : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GT2_GTXRXN_IN                           : in   std_logic;
    GT2_GTXRXP_IN                           : in   std_logic;
    GT2_RXCDRLOCK_OUT                       : out  std_logic;
    GT2_RXELECIDLE_OUT                      : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GT2_RXBUFRESET_IN                       : in   std_logic;
    GT2_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GT2_RXRESETDONE_OUT                     : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    GT2_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
    GT2_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);    
    GT2_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT2_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    GT2_TXDLYEN_IN                          : in   std_logic;
    GT2_TXDLYSRESET_IN                      : in   std_logic;
    GT2_TXDLYSRESETDONE_OUT                 : out  std_logic;
    GT2_TXPHALIGN_IN                        : in   std_logic;
    GT2_TXPHALIGNDONE_OUT                   : out  std_logic;
    GT2_TXPHALIGNEN_IN                      : in   std_logic;
    GT2_TXPHDLYRESET_IN                     : in   std_logic;
    GT2_TXPHINIT_IN                         : in   std_logic;
    GT2_TXPHINITDONE_OUT                    : out  std_logic;    
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT2_GTTXRESET_IN                        : in   std_logic;
    GT2_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    GT2_TXOUTCLK_OUT                        : out  std_logic;
    GT2_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT2_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT2_TXPCSRESET_IN                       : in   std_logic;
    GT2_TXUSRCLK_IN                         : in   std_logic;
    GT2_TXUSRCLK2_IN                        : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT2_GTXTXN_OUT                          : out  std_logic;
    GT2_GTXTXP_OUT                          : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GT2_TXRESETDONE_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GT2_TXPRBSFORCEERR_IN                   : in   std_logic;
    GT2_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GT2_TXELECIDLE_IN                       : in   std_logic;

    --GT3  (X0Y15)
    --____________________________CHANNEL PORTS________________________________
    ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
    GT3_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT3_DRPCLK_IN                           : in   std_logic;
    GT3_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT3_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT3_DRPEN_IN                            : in   std_logic;
    GT3_DRPRDY_OUT                          : out  std_logic;
    GT3_DRPWE_IN                            : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    GT3_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    GT3_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    GT3_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT3_TXPD_IN                             : in   std_logic_vector(1 downto 0);        
    ------------------------------- Receive Ports ------------------------------
    GT3_RXUSERRDY_IN                        : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GT3_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT3_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT3_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT3_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GT3_RXCHANBONDSEQ_OUT                   : out  std_logic;
    GT3_RXCHBONDEN_IN                       : in   std_logic;
    GT3_RXCHBONDI_IN                        : in   std_logic_vector(4 downto 0);
    GT3_RXCHBONDLEVEL_IN                    : in   std_logic_vector(2 downto 0);
    GT3_RXCHBONDMASTER_IN                   : in   std_logic;
    GT3_RXCHBONDO_OUT                       : out  std_logic_vector(4 downto 0);
    GT3_RXCHBONDSLAVE_IN                    : in   std_logic;
    ------------------- Receive Ports - Channel Bonding Ports  -----------------
    GT3_RXCHANISALIGNED_OUT                 : out  std_logic;
    GT3_RXCHANREALIGN_OUT                   : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GT3_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GT3_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT3_RXBYTEREALIGN_OUT                   : out  std_logic;
    GT3_RXCOMMADET_OUT                      : out  std_logic;
    GT3_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT3_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GT3_RXPRBSCNTRESET_IN                   : in   std_logic;
    GT3_RXPRBSERR_OUT                       : out  std_logic;
    GT3_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - RX Data Path interface -----------------
    GT3_GTRXRESET_IN                        : in   std_logic;
    GT3_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT3_RXOUTCLK_OUT                        : out  std_logic;    
    GT3_RXPCSRESET_IN                       : in   std_logic;
    GT3_RXUSRCLK_IN                         : in   std_logic;
    GT3_RXUSRCLK2_IN                        : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GT3_GTXRXN_IN                           : in   std_logic;
    GT3_GTXRXP_IN                           : in   std_logic;
    GT3_RXCDRLOCK_OUT                       : out  std_logic;
    GT3_RXELECIDLE_OUT                      : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GT3_RXBUFRESET_IN                       : in   std_logic;
    GT3_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GT3_RXRESETDONE_OUT                     : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    GT3_TXPOSTCURSOR_IN                     : in   std_logic_vector(4 downto 0);
    GT3_TXPRECURSOR_IN                      : in   std_logic_vector(4 downto 0);    
    GT3_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT3_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    GT3_TXDLYEN_IN                          : in   std_logic;
    GT3_TXDLYSRESET_IN                      : in   std_logic;
    GT3_TXDLYSRESETDONE_OUT                 : out  std_logic;
    GT3_TXPHALIGN_IN                        : in   std_logic;
    GT3_TXPHALIGNDONE_OUT                   : out  std_logic;
    GT3_TXPHALIGNEN_IN                      : in   std_logic;
    GT3_TXPHDLYRESET_IN                     : in   std_logic;
    GT3_TXPHINIT_IN                         : in   std_logic;
    GT3_TXPHINITDONE_OUT                    : out  std_logic;    
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT3_GTTXRESET_IN                        : in   std_logic;
    GT3_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    GT3_TXOUTCLK_OUT                        : out  std_logic;
    GT3_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT3_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT3_TXPCSRESET_IN                       : in   std_logic;
    GT3_TXUSRCLK_IN                         : in   std_logic;
    GT3_TXUSRCLK2_IN                        : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT3_GTXTXN_OUT                          : out  std_logic;
    GT3_GTXTXP_OUT                          : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GT3_TXRESETDONE_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GT3_TXPRBSFORCEERR_IN                   : in   std_logic;
    GT3_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GT3_TXELECIDLE_IN                       : in   std_logic;


    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT0_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT0_QPLLLOCK_OUT                        : out  std_logic;
    GT0_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_QPLLREFCLKLOST_OUT                  : out  std_logic;	
    GT0_QPLLRESET_IN                        : in   std_logic


);


end zynq_xaui_gt_wrapper;
    
architecture RTL of zynq_xaui_gt_wrapper is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "xaui_gt_wrapper,gtwizard_v2_2,{protocol_file=xaui}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;
    signal   gt0_qplloutclk_i         :   std_logic;
    signal   gt0_qplloutrefclk_i      :   std_logic;

  
    signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
    signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
  
 
    signal   gt0_qpllclk_i            :   std_logic;
    signal   gt0_qpllrefclk_i         :   std_logic;

    signal   gt1_qpllclk_i            :   std_logic;
    signal   gt1_qpllrefclk_i         :   std_logic;

    signal   gt2_qpllclk_i            :   std_logic;
    signal   gt2_qpllrefclk_i         :   std_logic;

    signal   gt3_qpllclk_i            :   std_logic;
    signal   gt3_qpllrefclk_i         :   std_logic;



--*************************** Component Declarations **************************
component zynq_xaui_gt_wrapper_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP       : string   := "false";
    RX_DFE_KL_CFG2_IN            : bit_vector :=   X"3010D90C";
    PMA_RSV_IN                   : bit_vector :=   X"00000000";
    PCS_RSVD_ATTR_IN             : bit_vector :=   X"000000000000";
    SIM_VERSION                  : string     := "4.0"

);
port 
(   
    ---------------------------------- Channel ---------------------------------
    QPLLCLK_IN                              : in   std_logic;
    QPLLREFCLK_IN                           : in   std_logic;
    ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
    DRPADDR_IN                              : in   std_logic_vector(8 downto 0);
    DRPCLK_IN                               : in   std_logic;
    DRPDI_IN                                : in   std_logic_vector(15 downto 0);
    DRPDO_OUT                               : out  std_logic_vector(15 downto 0);
    DRPEN_IN                                : in   std_logic;
    DRPRDY_OUT                              : out  std_logic;
    DRPWE_IN                                : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    EYESCANDATAERROR_OUT                    : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    LOOPBACK_IN                             : in   std_logic_vector(2 downto 0);
    RXPD_IN                                 : in   std_logic_vector(1 downto 0);
    TXPD_IN                                 : in   std_logic_vector(1 downto 0);        
    ------------------------------- Receive Ports ------------------------------
    RXUSERRDY_IN                            : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    RXCHARISCOMMA_OUT                       : out  std_logic_vector(1 downto 0);
    RXCHARISK_OUT                           : out  std_logic_vector(1 downto 0);
    RXDISPERR_OUT                           : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE_OUT                        : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    RXCHANBONDSEQ_OUT                       : out  std_logic;
    RXCHBONDEN_IN                           : in   std_logic;
    RXCHBONDI_IN                            : in   std_logic_vector(4 downto 0);
    RXCHBONDLEVEL_IN                        : in   std_logic_vector(2 downto 0);
    RXCHBONDMASTER_IN                       : in   std_logic;
    RXCHBONDO_OUT                           : out  std_logic_vector(4 downto 0);
    RXCHBONDSLAVE_IN                        : in   std_logic;
    ------------------- Receive Ports - Channel Bonding Ports  -----------------
    RXCHANISALIGNED_OUT                     : out  std_logic;
    RXCHANREALIGN_OUT                       : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    RXCLKCORCNT_OUT                         : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    RXBYTEISALIGNED_OUT                     : out  std_logic;
    RXBYTEREALIGN_OUT                       : out  std_logic;
    RXCOMMADET_OUT                          : out  std_logic;
    RXMCOMMAALIGNEN_IN                      : in   std_logic;
    RXPCOMMAALIGNEN_IN                      : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    RXPRBSCNTRESET_IN                       : in   std_logic;
    RXPRBSERR_OUT                           : out  std_logic;
    RXPRBSSEL_IN                            : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - RX Data Path interface -----------------
    GTRXRESET_IN                            : in   std_logic;
    RXDATA_OUT                              : out  std_logic_vector(15 downto 0);
    RXOUTCLK_OUT                            : out  std_logic;    
    RXPCSRESET_IN                           : in   std_logic;
    RXUSRCLK_IN                             : in   std_logic;
    RXUSRCLK2_IN                            : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTXRXN_IN                               : in   std_logic;
    GTXRXP_IN                               : in   std_logic;
    RXCDRLOCK_OUT                           : out  std_logic;
    RXELECIDLE_OUT                          : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    RXBUFRESET_IN                           : in   std_logic;
    RXBUFSTATUS_OUT                         : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    RXRESETDONE_OUT                         : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    TXPOSTCURSOR_IN                         : in   std_logic_vector(4 downto 0);
    TXPRECURSOR_IN                          : in   std_logic_vector(4 downto 0);    
    TXUSERRDY_IN                            : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TXCHARISK_IN                            : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    TXDLYEN_IN                              : in   std_logic;
    TXDLYSRESET_IN                          : in   std_logic;
    TXDLYSRESETDONE_OUT                     : out  std_logic;
    TXPHALIGN_IN                            : in   std_logic;
    TXPHALIGNDONE_OUT                       : out  std_logic;
    TXPHALIGNEN_IN                          : in   std_logic;
    TXPHDLYRESET_IN                         : in   std_logic;
    TXPHINIT_IN                             : in   std_logic;
    TXPHINITDONE_OUT                        : out  std_logic;    
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTTXRESET_IN                            : in   std_logic;
    TXDATA_IN                               : in   std_logic_vector(15 downto 0);
    TXOUTCLK_OUT                            : out  std_logic;
    TXOUTCLKFABRIC_OUT                      : out  std_logic;
    TXOUTCLKPCS_OUT                         : out  std_logic;
    TXPCSRESET_IN                           : in   std_logic;
    TXUSRCLK_IN                             : in   std_logic;
    TXUSRCLK2_IN                            : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTXTXN_OUT                              : out  std_logic;
    GTXTXP_OUT                              : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    TXRESETDONE_OUT                         : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    TXPRBSFORCEERR_IN                       : in   std_logic;
    TXPRBSSEL_IN                            : in   std_logic_vector(2 downto 0);
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    TXELECIDLE_IN                           : in   std_logic


);
end component;



--*************************Logic to set Attribute QPLL_FB_DIV*****************************
    impure function conv_qpll_fbdiv_top (qpllfbdiv_top : in integer) return bit_vector is
    begin
       if (qpllfbdiv_top = 16) then
         return "0000100000";
       elsif (qpllfbdiv_top = 20) then
         return "0000110000" ;
       elsif (qpllfbdiv_top = 32) then
         return "0001100000" ;
       elsif (qpllfbdiv_top = 40) then
         return "0010000000" ;
       elsif (qpllfbdiv_top = 64) then
         return "0011100000" ;
       elsif (qpllfbdiv_top = 66) then
         return "0101000000" ;
       elsif (qpllfbdiv_top = 80) then
         return "0100100000" ;
       elsif (qpllfbdiv_top = 100) then
         return "0101110000" ;
       else 
         return "0000000000" ;
       end if;
    end function;

    impure function conv_qpll_fbdiv_ratio (qpllfbdiv_top : in integer) return bit is
    begin
       if (qpllfbdiv_top = 16) then
         return '1';
       elsif (qpllfbdiv_top = 20) then
         return '1' ;
       elsif (qpllfbdiv_top = 32) then
         return '1' ;
       elsif (qpllfbdiv_top = 40) then
         return '1' ;
       elsif (qpllfbdiv_top = 64) then
         return '1' ;
       elsif (qpllfbdiv_top = 66) then
         return '0' ;
       elsif (qpllfbdiv_top = 80) then
         return '1' ;
       elsif (qpllfbdiv_top = 100) then
         return '1' ;
       else 
         return '1' ;
       end if;
    end function;

    constant   QPLL_FBDIV_IN    :   bit_vector(9 downto 0) := conv_qpll_fbdiv_top(QPLL_FBDIV_TOP);
    constant   QPLL_FBDIV_RATIO :   bit := conv_qpll_fbdiv_ratio(QPLL_FBDIV_TOP);

--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';

    gt0_qpllclk_i    <= gt0_qplloutclk_i;  
    gt0_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt1_qpllclk_i    <= gt0_qplloutclk_i;  
    gt1_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt2_qpllclk_i    <= gt0_qplloutclk_i;  
    gt2_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    gt3_qpllclk_i    <= gt0_qplloutclk_i;  
    gt3_qpllrefclk_i <= gt0_qplloutrefclk_i; 

    --------------------------- GT Instances  -------------------------------   

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y12)

    gt0_zynq_xaui_gt_wrapper_i : zynq_xaui_gt_wrapper_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000002",
        SIM_VERSION                   =>  SIM_VERSION  
        
    )
    port map
    (
        ---------------------------------- Channel ---------------------------------
        QPLLCLK_IN                      =>      gt0_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt0_qpllrefclk_i,
        ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
        DRPADDR_IN                      =>      GT0_DRPADDR_IN,
        DRPCLK_IN                       =>      GT0_DRPCLK_IN,
        DRPDI_IN                        =>      GT0_DRPDI_IN,
        DRPDO_OUT                       =>      GT0_DRPDO_OUT,
        DRPEN_IN                        =>      GT0_DRPEN_IN,
        DRPRDY_OUT                      =>      GT0_DRPRDY_OUT,
        DRPWE_IN                        =>      GT0_DRPWE_IN,
        ------------------------------- Eye Scan Ports -----------------------------
        EYESCANDATAERROR_OUT            =>      GT0_EYESCANDATAERROR_OUT,
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GT0_LOOPBACK_IN,
        RXPD_IN                         =>      GT0_RXPD_IN,
        TXPD_IN                         =>      GT0_TXPD_IN,        
        ------------------------------- Receive Ports ------------------------------
        RXUSERRDY_IN                    =>      GT0_RXUSERRDY_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GT0_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT0_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GT0_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT0_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GT0_RXCHANBONDSEQ_OUT,
        RXCHBONDEN_IN                   =>      GT0_RXCHBONDEN_IN,
        RXCHBONDI_IN                    =>      GT0_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GT0_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GT0_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GT0_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GT0_RXCHBONDSLAVE_IN,
        ------------------- Receive Ports - Channel Bonding Ports  -----------------
        RXCHANISALIGNED_OUT             =>      GT0_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GT0_RXCHANREALIGN_OUT,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GT0_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GT0_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT0_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT0_RXCOMMADET_OUT,
        RXMCOMMAALIGNEN_IN              =>      GT0_RXMCOMMAALIGNEN_IN,
        RXPCOMMAALIGNEN_IN              =>      GT0_RXPCOMMAALIGNEN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        RXPRBSCNTRESET_IN               =>      GT0_RXPRBSCNTRESET_IN,
        RXPRBSERR_OUT                   =>      GT0_RXPRBSERR_OUT,
        RXPRBSSEL_IN                    =>      GT0_RXPRBSSEL_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        GTRXRESET_IN                    =>      GT0_GTRXRESET_IN,
        RXDATA_OUT                      =>      GT0_RXDATA_OUT,
        RXOUTCLK_OUT                    =>      GT0_RXOUTCLK_OUT,        
        RXPCSRESET_IN                   =>      GT0_RXPCSRESET_IN,
        RXUSRCLK_IN                     =>      GT0_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT0_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        GTXRXN_IN                       =>      GT0_GTXRXN_IN,
        GTXRXP_IN                       =>      GT0_GTXRXP_IN,
        RXCDRLOCK_OUT                   =>      GT0_RXCDRLOCK_OUT,
        RXELECIDLE_OUT                  =>      GT0_RXELECIDLE_OUT,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GT0_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GT0_RXBUFSTATUS_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        RXRESETDONE_OUT                 =>      GT0_RXRESETDONE_OUT,
        ------------------------------- Transmit Ports -----------------------------
        TXPOSTCURSOR_IN                 =>      GT0_TXPOSTCURSOR_IN,
        TXPRECURSOR_IN                  =>      GT0_TXPRECURSOR_IN,
        TXUSERRDY_IN                    =>      GT0_TXUSERRDY_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GT0_TXCHARISK_IN,
        ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
        TXDLYEN_IN                      =>      GT0_TXDLYEN_IN,
        TXDLYSRESET_IN                  =>      GT0_TXDLYSRESET_IN,
        TXDLYSRESETDONE_OUT             =>      GT0_TXDLYSRESETDONE_OUT,
        TXPHALIGN_IN                    =>      GT0_TXPHALIGN_IN,
        TXPHALIGNDONE_OUT               =>      GT0_TXPHALIGNDONE_OUT,
        TXPHALIGNEN_IN                  =>      GT0_TXPHALIGNEN_IN,
        TXPHDLYRESET_IN                 =>      GT0_TXPHDLYRESET_IN,
        TXPHINIT_IN                     =>      GT0_TXPHINIT_IN,
        TXPHINITDONE_OUT                =>      GT0_TXPHINITDONE_OUT,        
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GTTXRESET_IN                    =>      GT0_GTTXRESET_IN,
        TXDATA_IN                       =>      GT0_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GT0_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT0_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT0_TXOUTCLKPCS_OUT,
        TXPCSRESET_IN                   =>      GT0_TXPCSRESET_IN,
        TXUSRCLK_IN                     =>      GT0_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT0_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT0_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT0_GTXTXP_OUT,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        TXRESETDONE_OUT                 =>      GT0_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXPRBSFORCEERR_IN               =>      GT0_TXPRBSFORCEERR_IN,
        TXPRBSSEL_IN                    =>      GT0_TXPRBSSEL_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GT0_TXELECIDLE_IN

    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y13)

    gt1_zynq_xaui_gt_wrapper_i : zynq_xaui_gt_wrapper_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000002",
        SIM_VERSION                   =>  SIM_VERSION 
        
    )
    port map
    (
        ---------------------------------- Channel ---------------------------------
        QPLLCLK_IN                      =>      gt1_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt1_qpllrefclk_i,
        ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
        DRPADDR_IN                      =>      GT1_DRPADDR_IN,
        DRPCLK_IN                       =>      GT1_DRPCLK_IN,
        DRPDI_IN                        =>      GT1_DRPDI_IN,
        DRPDO_OUT                       =>      GT1_DRPDO_OUT,
        DRPEN_IN                        =>      GT1_DRPEN_IN,
        DRPRDY_OUT                      =>      GT1_DRPRDY_OUT,
        DRPWE_IN                        =>      GT1_DRPWE_IN,
        ------------------------------- Eye Scan Ports -----------------------------
        EYESCANDATAERROR_OUT            =>      GT1_EYESCANDATAERROR_OUT,
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GT1_LOOPBACK_IN,
        RXPD_IN                         =>      GT1_RXPD_IN,
        TXPD_IN                         =>      GT1_TXPD_IN,        
        ------------------------------- Receive Ports ------------------------------
        RXUSERRDY_IN                    =>      GT1_RXUSERRDY_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GT1_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT1_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GT1_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT1_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GT1_RXCHANBONDSEQ_OUT,
        RXCHBONDEN_IN                   =>      GT1_RXCHBONDEN_IN,
        RXCHBONDI_IN                    =>      GT1_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GT1_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GT1_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GT1_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GT1_RXCHBONDSLAVE_IN,
        ------------------- Receive Ports - Channel Bonding Ports  -----------------
        RXCHANISALIGNED_OUT             =>      GT1_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GT1_RXCHANREALIGN_OUT,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GT1_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GT1_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT1_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT1_RXCOMMADET_OUT,
        RXMCOMMAALIGNEN_IN              =>      GT1_RXMCOMMAALIGNEN_IN,
        RXPCOMMAALIGNEN_IN              =>      GT1_RXPCOMMAALIGNEN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        RXPRBSCNTRESET_IN               =>      GT1_RXPRBSCNTRESET_IN,
        RXPRBSERR_OUT                   =>      GT1_RXPRBSERR_OUT,
        RXPRBSSEL_IN                    =>      GT1_RXPRBSSEL_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        GTRXRESET_IN                    =>      GT1_GTRXRESET_IN,
        RXDATA_OUT                      =>      GT1_RXDATA_OUT,
        RXOUTCLK_OUT                    =>      GT1_RXOUTCLK_OUT,        
        RXPCSRESET_IN                   =>      GT1_RXPCSRESET_IN,
        RXUSRCLK_IN                     =>      GT1_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT1_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        GTXRXN_IN                       =>      GT1_GTXRXN_IN,
        GTXRXP_IN                       =>      GT1_GTXRXP_IN,
        RXCDRLOCK_OUT                   =>      GT1_RXCDRLOCK_OUT,
        RXELECIDLE_OUT                  =>      GT1_RXELECIDLE_OUT,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GT1_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GT1_RXBUFSTATUS_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        RXRESETDONE_OUT                 =>      GT1_RXRESETDONE_OUT,
        ------------------------------- Transmit Ports -----------------------------
        TXPOSTCURSOR_IN                 =>      GT1_TXPOSTCURSOR_IN,
        TXPRECURSOR_IN                  =>      GT1_TXPRECURSOR_IN,
        TXUSERRDY_IN                    =>      GT1_TXUSERRDY_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GT1_TXCHARISK_IN,
        ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
        TXDLYEN_IN                      =>      GT1_TXDLYEN_IN,
        TXDLYSRESET_IN                  =>      GT1_TXDLYSRESET_IN,
        TXDLYSRESETDONE_OUT             =>      GT1_TXDLYSRESETDONE_OUT,
        TXPHALIGN_IN                    =>      GT1_TXPHALIGN_IN,
        TXPHALIGNDONE_OUT               =>      GT1_TXPHALIGNDONE_OUT,
        TXPHALIGNEN_IN                  =>      GT1_TXPHALIGNEN_IN,
        TXPHDLYRESET_IN                 =>      GT1_TXPHDLYRESET_IN,
        TXPHINIT_IN                     =>      GT1_TXPHINIT_IN,
        TXPHINITDONE_OUT                =>      GT1_TXPHINITDONE_OUT,        
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GTTXRESET_IN                    =>      GT1_GTTXRESET_IN,
        TXDATA_IN                       =>      GT1_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GT1_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT1_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT1_TXOUTCLKPCS_OUT,
        TXPCSRESET_IN                   =>      GT1_TXPCSRESET_IN,
        TXUSRCLK_IN                     =>      GT1_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT1_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT1_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT1_GTXTXP_OUT,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        TXRESETDONE_OUT                 =>      GT1_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXPRBSFORCEERR_IN               =>      GT1_TXPRBSFORCEERR_IN,
        TXPRBSSEL_IN                    =>      GT1_TXPRBSSEL_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GT1_TXELECIDLE_IN

    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y14)

    gt2_zynq_xaui_gt_wrapper_i : zynq_xaui_gt_wrapper_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000002",
        SIM_VERSION                   =>  SIM_VERSION    
        
    )
    port map
    (
        ---------------------------------- Channel ---------------------------------
        QPLLCLK_IN                      =>      gt2_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt2_qpllrefclk_i,
        ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
        DRPADDR_IN                      =>      GT2_DRPADDR_IN,
        DRPCLK_IN                       =>      GT2_DRPCLK_IN,
        DRPDI_IN                        =>      GT2_DRPDI_IN,
        DRPDO_OUT                       =>      GT2_DRPDO_OUT,
        DRPEN_IN                        =>      GT2_DRPEN_IN,
        DRPRDY_OUT                      =>      GT2_DRPRDY_OUT,
        DRPWE_IN                        =>      GT2_DRPWE_IN,
        ------------------------------- Eye Scan Ports -----------------------------
        EYESCANDATAERROR_OUT            =>      GT2_EYESCANDATAERROR_OUT,
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GT2_LOOPBACK_IN,
        RXPD_IN                         =>      GT2_RXPD_IN,
        TXPD_IN                         =>      GT2_TXPD_IN,        
        ------------------------------- Receive Ports ------------------------------
        RXUSERRDY_IN                    =>      GT2_RXUSERRDY_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GT2_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT2_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GT2_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT2_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GT2_RXCHANBONDSEQ_OUT,
        RXCHBONDEN_IN                   =>      GT2_RXCHBONDEN_IN,
        RXCHBONDI_IN                    =>      GT2_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GT2_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GT2_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GT2_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GT2_RXCHBONDSLAVE_IN,
        ------------------- Receive Ports - Channel Bonding Ports  -----------------
        RXCHANISALIGNED_OUT             =>      GT2_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GT2_RXCHANREALIGN_OUT,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GT2_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GT2_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT2_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT2_RXCOMMADET_OUT,
        RXMCOMMAALIGNEN_IN              =>      GT2_RXMCOMMAALIGNEN_IN,
        RXPCOMMAALIGNEN_IN              =>      GT2_RXPCOMMAALIGNEN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        RXPRBSCNTRESET_IN               =>      GT2_RXPRBSCNTRESET_IN,
        RXPRBSERR_OUT                   =>      GT2_RXPRBSERR_OUT,
        RXPRBSSEL_IN                    =>      GT2_RXPRBSSEL_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        GTRXRESET_IN                    =>      GT2_GTRXRESET_IN,
        RXDATA_OUT                      =>      GT2_RXDATA_OUT,
        RXOUTCLK_OUT                    =>      GT2_RXOUTCLK_OUT,        
        RXPCSRESET_IN                   =>      GT2_RXPCSRESET_IN,
        RXUSRCLK_IN                     =>      GT2_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT2_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        GTXRXN_IN                       =>      GT2_GTXRXN_IN,
        GTXRXP_IN                       =>      GT2_GTXRXP_IN,
        RXCDRLOCK_OUT                   =>      GT2_RXCDRLOCK_OUT,
        RXELECIDLE_OUT                  =>      GT2_RXELECIDLE_OUT,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GT2_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GT2_RXBUFSTATUS_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        RXRESETDONE_OUT                 =>      GT2_RXRESETDONE_OUT,
        ------------------------------- Transmit Ports -----------------------------
        TXPOSTCURSOR_IN                 =>      GT2_TXPOSTCURSOR_IN,
        TXPRECURSOR_IN                  =>      GT2_TXPRECURSOR_IN,
        TXUSERRDY_IN                    =>      GT2_TXUSERRDY_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GT2_TXCHARISK_IN,
        ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
        TXDLYEN_IN                      =>      GT2_TXDLYEN_IN,
        TXDLYSRESET_IN                  =>      GT2_TXDLYSRESET_IN,
        TXDLYSRESETDONE_OUT             =>      GT2_TXDLYSRESETDONE_OUT,
        TXPHALIGN_IN                    =>      GT2_TXPHALIGN_IN,
        TXPHALIGNDONE_OUT               =>      GT2_TXPHALIGNDONE_OUT,
        TXPHALIGNEN_IN                  =>      GT2_TXPHALIGNEN_IN,
        TXPHDLYRESET_IN                 =>      GT2_TXPHDLYRESET_IN,
        TXPHINIT_IN                     =>      GT2_TXPHINIT_IN,
        TXPHINITDONE_OUT                =>      GT2_TXPHINITDONE_OUT,        
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GTTXRESET_IN                    =>      GT2_GTTXRESET_IN,
        TXDATA_IN                       =>      GT2_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GT2_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT2_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT2_TXOUTCLKPCS_OUT,
        TXPCSRESET_IN                   =>      GT2_TXPCSRESET_IN,
        TXUSRCLK_IN                     =>      GT2_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT2_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT2_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT2_GTXTXP_OUT,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        TXRESETDONE_OUT                 =>      GT2_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXPRBSFORCEERR_IN               =>      GT2_TXPRBSFORCEERR_IN,
        TXPRBSSEL_IN                    =>      GT2_TXPRBSSEL_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GT2_TXELECIDLE_IN

    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y15)

    gt3_zynq_xaui_gt_wrapper_i : zynq_xaui_gt_wrapper_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP        =>  WRAPPER_SIM_GTRESET_SPEEDUP,
        RX_DFE_KL_CFG2_IN             =>  RX_DFE_KL_CFG2_IN,
        PMA_RSV_IN                    =>  PMA_RSV_IN,
        PCS_RSVD_ATTR_IN              =>  X"000000000002",
        SIM_VERSION                   =>  SIM_VERSION
        
    )
    port map
    (
        ---------------------------------- Channel ---------------------------------
        QPLLCLK_IN                      =>      gt3_qpllclk_i,
        QPLLREFCLK_IN                   =>      gt3_qpllrefclk_i,
        ---------------- Channel - Dynamic Reconfiguration Port (DRP) --------------
        DRPADDR_IN                      =>      GT3_DRPADDR_IN,
        DRPCLK_IN                       =>      GT3_DRPCLK_IN,
        DRPDI_IN                        =>      GT3_DRPDI_IN,
        DRPDO_OUT                       =>      GT3_DRPDO_OUT,
        DRPEN_IN                        =>      GT3_DRPEN_IN,
        DRPRDY_OUT                      =>      GT3_DRPRDY_OUT,
        DRPWE_IN                        =>      GT3_DRPWE_IN,
        ------------------------------- Eye Scan Ports -----------------------------
        EYESCANDATAERROR_OUT            =>      GT3_EYESCANDATAERROR_OUT,
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GT3_LOOPBACK_IN,
        RXPD_IN                         =>      GT3_RXPD_IN,
        TXPD_IN                         =>      GT3_TXPD_IN,        
        ------------------------------- Receive Ports ------------------------------
        RXUSERRDY_IN                    =>      GT3_RXUSERRDY_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GT3_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GT3_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GT3_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GT3_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GT3_RXCHANBONDSEQ_OUT,
        RXCHBONDEN_IN                   =>      GT3_RXCHBONDEN_IN,
        RXCHBONDI_IN                    =>      GT3_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GT3_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GT3_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GT3_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GT3_RXCHBONDSLAVE_IN,
        ------------------- Receive Ports - Channel Bonding Ports  -----------------
        RXCHANISALIGNED_OUT             =>      GT3_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GT3_RXCHANREALIGN_OUT,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GT3_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GT3_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GT3_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GT3_RXCOMMADET_OUT,
        RXMCOMMAALIGNEN_IN              =>      GT3_RXMCOMMAALIGNEN_IN,
        RXPCOMMAALIGNEN_IN              =>      GT3_RXPCOMMAALIGNEN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        RXPRBSCNTRESET_IN               =>      GT3_RXPRBSCNTRESET_IN,
        RXPRBSERR_OUT                   =>      GT3_RXPRBSERR_OUT,
        RXPRBSSEL_IN                    =>      GT3_RXPRBSSEL_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        GTRXRESET_IN                    =>      GT3_GTRXRESET_IN,
        RXDATA_OUT                      =>      GT3_RXDATA_OUT,
        RXOUTCLK_OUT                    =>      GT3_RXOUTCLK_OUT,        
        RXPCSRESET_IN                   =>      GT3_RXPCSRESET_IN,
        RXUSRCLK_IN                     =>      GT3_RXUSRCLK_IN,
        RXUSRCLK2_IN                    =>      GT3_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        GTXRXN_IN                       =>      GT3_GTXRXN_IN,
        GTXRXP_IN                       =>      GT3_GTXRXP_IN,
        RXCDRLOCK_OUT                   =>      GT3_RXCDRLOCK_OUT,
        RXELECIDLE_OUT                  =>      GT3_RXELECIDLE_OUT,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GT3_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GT3_RXBUFSTATUS_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        RXRESETDONE_OUT                 =>      GT3_RXRESETDONE_OUT,
        ------------------------------- Transmit Ports -----------------------------
        TXPOSTCURSOR_IN                 =>      GT3_TXPOSTCURSOR_IN,
        TXPRECURSOR_IN                  =>      GT3_TXPRECURSOR_IN,
        TXUSERRDY_IN                    =>      GT3_TXUSERRDY_IN,        
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GT3_TXCHARISK_IN,
        ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
        TXDLYEN_IN                      =>      GT3_TXDLYEN_IN,
        TXDLYSRESET_IN                  =>      GT3_TXDLYSRESET_IN,
        TXDLYSRESETDONE_OUT             =>      GT3_TXDLYSRESETDONE_OUT,
        TXPHALIGN_IN                    =>      GT3_TXPHALIGN_IN,
        TXPHALIGNDONE_OUT               =>      GT3_TXPHALIGNDONE_OUT,
        TXPHALIGNEN_IN                  =>      GT3_TXPHALIGNEN_IN,
        TXPHDLYRESET_IN                 =>      GT3_TXPHDLYRESET_IN,
        TXPHINIT_IN                     =>      GT3_TXPHINIT_IN,
        TXPHINITDONE_OUT                =>      GT3_TXPHINITDONE_OUT,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GTTXRESET_IN                    =>      GT3_GTTXRESET_IN,
        TXDATA_IN                       =>      GT3_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GT3_TXOUTCLK_OUT,
        TXOUTCLKFABRIC_OUT              =>      GT3_TXOUTCLKFABRIC_OUT,
        TXOUTCLKPCS_OUT                 =>      GT3_TXOUTCLKPCS_OUT,
        TXPCSRESET_IN                   =>      GT3_TXPCSRESET_IN,
        TXUSRCLK_IN                     =>      GT3_TXUSRCLK_IN,
        TXUSRCLK2_IN                    =>      GT3_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTXTXN_OUT                      =>      GT3_GTXTXN_OUT,
        GTXTXP_OUT                      =>      GT3_GTXTXP_OUT,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        TXRESETDONE_OUT                 =>      GT3_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXPRBSFORCEERR_IN               =>      GT3_TXPRBSFORCEERR_IN,
        TXPRBSSEL_IN                    =>      GT3_TXPRBSSEL_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GT3_TXELECIDLE_IN

    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTXE2_COMMON____________________________________

    gtxe2_common_0_i : GTXE2_COMMON
    generic map
    (
            -- Simulation attributes
            SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
            SIM_QPLLREFCLK_SEL   => ("001"),
            SIM_VERSION          => SIM_VERSION,


       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000040000001000"),
        COMMON_CFG                              =>     (x"00000000"),
        QPLL_CFG                                =>     (x"06801C1"),
        QPLL_CLKOUT_CFG                         =>     ("0000"),
        QPLL_COARSE_FREQ_OVRD                   =>     ("010000"),
        QPLL_COARSE_FREQ_OVRD_EN                =>     ('0'),
        QPLL_CP                                 =>     ("0000011111"),
        QPLL_CP_MONITOR_EN                      =>     ('0'),
        QPLL_DMONITOR_SEL                       =>     ('0'),
        QPLL_FBDIV                              =>     (QPLL_FBDIV_IN),
        QPLL_FBDIV_MONITOR_EN                   =>     ('0'),
        QPLL_FBDIV_RATIO                        =>     (QPLL_FBDIV_RATIO),
        QPLL_INIT_CFG                           =>     (x"000006"),
        QPLL_LOCK_CFG                           =>     (x"21E8"),
        QPLL_LPF                                =>     ("1111"),
        QPLL_REFCLK_DIV                         =>     (1)

        
    )
    port map
    (
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      tied_to_ground_vec_i(7 downto 0),
        DRPCLK                          =>      tied_to_ground_i,
        DRPDI                           =>      tied_to_ground_vec_i(15 downto 0),
        DRPDO                           =>      open,
        DRPEN                           =>      tied_to_ground_i,
        DRPRDY                          =>      open,
        DRPWE                           =>      tied_to_ground_i,
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GTGREFCLK                       =>      tied_to_ground_i,
        GTNORTHREFCLK0                  =>      tied_to_ground_i,
        GTNORTHREFCLK1                  =>      tied_to_ground_i,
        GTREFCLK0                       =>      GT0_GTREFCLK0_COMMON_IN,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTSOUTHREFCLK0                  =>      tied_to_ground_i,
        GTSOUTHREFCLK1                  =>      tied_to_ground_i,
        ------------------------- Common Block - QPLL Ports ------------------------
        QPLLDMONITOR                    =>      open,		
        QPLLFBCLKLOST                   =>      open,
        QPLLLOCK                        =>      GT0_QPLLLOCK_OUT,
        QPLLLOCKDETCLK                  =>      GT0_QPLLLOCKDETCLK_IN,
        QPLLLOCKEN                      =>      tied_to_vcc_i,
        QPLLOUTCLK                      =>      gt0_qplloutclk_i,
        QPLLOUTREFCLK                   =>      gt0_qplloutrefclk_i,
        QPLLOUTRESET                    =>      tied_to_ground_i,
        QPLLPD                          =>      tied_to_ground_i,
        QPLLREFCLKLOST                  =>      GT0_QPLLREFCLKLOST_OUT,
        QPLLREFCLKSEL                   =>      "001",
        QPLLRESET                       =>      GT0_QPLLRESET_IN,
        QPLLRSVD1                       =>      "0000000000000000",
        QPLLRSVD2                       =>      "11111",
        REFCLKOUTMONITOR                =>      open,
        ----------------------------- Common Block Ports ---------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i
    );

     
end RTL;
