XlxV64EB    9423    1890�bbA����/2�֪T����%�����=F�$<�cτ3���Z��+����m���R4����F�O����H����o�ZA9V��0`E����Q���Q��p[�>:N�� y�"o��(�YW���_���4��Ia,��v�i�7D���߸�mʞy#�_#P��0
��$�����dļ�������m�3��{#*b��<0�eZx瘜�ޯ��?<�!y���G8�LF��r��2�:��S���=^���R&f���M��ϗ�LD��i'�S�FYOIR�c�>G?��C@�.��Chi�a5G�eжJf$�-],㠎.��8\�y��,	�]�	�Q}��i�KS��(��;�"\T�d���/���<0C�-���0��BQ�+	v�l�Ho�7P���sM�a�M��b<g4	��s�B���f>*a�)���������Á���xyF#+���s'�fΘ��	/[�9��//"ɷ��q��\�)����o���n	��+
.
 ��y�
�s��.~q�fX<��O� ����NN{[��huG�ʸ��{�IW�q��@C'��� ��6'����@M����K� pԐ�}�w�K�����-!ާ�y��SЦ[����Cy�BJR�`d�<�N� �
R3��S|Q]�^3z|�)�3��p⟞P\�0�%h��;_��(=v����-Z�,j�������f0]�I���曧l�h#G��1�9�� ��I9ֱbE渻B��bN�.�F�xƹ���Xl�x���r�َ22	fYɉGG����ª��_�QG�k̓U�)A������%F�*���C��L��E���6���~r�6��#�=�����ԩ����6v��އ��CyH��م�7�x�{ȝ�a�  ��-����y���R���˵6 ��X�IՎוtƁU�ώף�!�'?C�&���U��&���}�2�j�T������b���m�=���{����&�y�WG���7m�aMtZ�& ��w�;���a0�:�M[Q���I3F�­�D�QL�3��Nl�\p�*1 dd�*���X��y�^�),�K�Y�����W�wz
��;�JR<�< ���h_��e�:�g�������6q�M���||$+G�(�S�!Զŝ�������m�ؠ�𧻓+��))?�
��_)�6؋�)��'�ü�oq�k�v�;3J�&�<��D����&��F�C�k�N�ʚ�MȨ0��j���s����\��11���O�|�l�kfu�]�Đ���
��S
��%C���=���)�A�{�m�ʩ+����^��v�T7�-�,��{B���.�{��k�#���%f� K!���L�`֚k�존v�Ia;��1��5jU���L�H��Z�bU�6�xy�����2����Y}[�E�YOd1_�j�>r���q��{�0e�6I�����47�V%�!t���^}���ϛ+[Фu��o�΄m�5c��N�?�~�ȈrrZ���`�o+�8����a�/���v&�	�tq�Z�jv� �;XJt��{c!��j�9��f�-���h�$���#2^����|RϸP.�u�b�5 y>�*�������늊�R�F�h�3 �t;�yE�R#�3Ooߨ��񑫡j9���(4�  D#�Cs�ht�-"���?x(�sS}�uN���f4uqw�'�H�AMJHʂ.pcݨ}�;^�y<��%fObS����T@ո���#f.��`)�[o�Q�"��K�9���|���`��b>LI���>ai��&�������N�ISi�*�W��Ý6������'�JhM�}q��v�p�Y�W	��������J��D�<��L�bD
�w����E�N���#�TPa9���1���/{���=u�M1jK��<7M@��e	�2eG@��`������c�Mm��7Zh�L����C�:{Mp�L����$3������DxhBz���C"�$�{��+���bV���jK�^��y�L��Վ�?���ҫ�Q�)��h��Y����)�z�d��c�6�~-ϻ��g�vKy�M���<.q�n��3X%�B���%h��j�N'��r��)��&�)1<����yt�o��P3�*�<�X>�F7�J��T5f��nݡ��<���Kz�Ƈjڎ�yNK�o򻽪��/��8T�B-Zr2|�+��D�i��}�c���)q�]�R�� <K�V�s���THR��U�c9JAx��+7�\]'$����P�a���֙����DZ��G}ڷBN�if���|�O���H���j�I<��D��ee�V��,G�3��L.�:��S��&��.��r�F��[�?�=��Y̷Ëj��%Qj"��0-�&�`Qp1\x`j2�����p�!n�`�غ���'�h�a��l%��R$�Di��Q��E�6��c��ΦzQ�HB��f5~�� �'���!{"�'"R���f��$�uy� ��kN���[�i*�����书c8A�<���^�1Xm�S��2vrAߤ����C+�-~j����M?��W���k��c̔ѻ�{B�cu$��Sb�w�����O�'1��ײ��C��/.�+�� Ⱥ�m��H��Ӿ>���ˍ������R�H�I�	t�\]SMV�$Q��H]X��l2���y/������a�Q���d���7#2�rK:W�T,#@�K���1)���+`.΂����,ջ��<M�j�~K8%I�b������|	-Ӯ��S��8���e�`p\��18[M�����_a[�=tJ��6o����*rb9'�:�̠b�����8��;`����%�� :�NU$/AZ�xv�9:�tC�`�.��X�.m2��QzA�n�0�"+���3p
�Ԣ/B}���X ��p*� ȢW�8WC1�0N��E������F)��=*wo��Hi�Ý�r5I9�Q��ぽk�w��O��H�(c�s��4[J	����?�a �?���9���$����0��-0�(�buQ/��EנeͲ����HsW�V���^m�[�'yIC�GSR؎�E�z8�te��p�H\@J�X��f2e��g�H��聐nܾ�Z�mr�T��|�k/����'�ӷ*4b�X��B���d���k��JM8��}���J�� ��G�e���@��'	C���E���S=VO0�d�{������4/��<��j��q0r�4�� �}����:��?l�y�w�2%p%'�_͂�su�\��8���,��d�)�{�����c��Wk�Swl�>�?�g�-��_�"jm���/��o��)�fcX���X�!�\'�����{SA3�'l�{��%JA�ף?�H�������.���s����BO�X�!w����-���>��Rh��ȹ`�X#�%��}�xznɝZ���B�%Y�X��*`y�z�"@£�ڛy�=.s���5���p�l�@'�O�ŕJhى.Ci���`���f�j���t��olU�e��hv����Â|ـ|�
9�K��EU���wQQ�ʾ����ˆY[!ȜΥEdhyȏ�l�a��C9�ݻr�n��34ME �`;��=�g��d��ޣ�ԛ����ɛ�D��`(-k;�n��/�(s�Ԑ��9��i�R�6@O�䭌Ֆ6�nf@��{�]�;3��$����[[ *;�f��4u���tI�\
 �!Ks#>h�Q+���{+-��6���X�]��ST��8�8ch�8U���`;���ۿ~%t�Yx��L��C��~���7�K.��d�*�7.�`�ҹ���uk��--3~R�-��l[E#���/�hg�p��ӽ�*�;�H9�����
�p�pO���Dh=��H8��p�6���G�����5�>Z�%)�2]�|�8_����\wy���8 ����F�1��t�kü&�P������N���:�s|�(Z�����=L�4Ԍa�y��.7��:�W�-�F��b�Z��$�U*�r1
��٠_��B�6��P��t�'�2��f�
Aa(Q-+���=������������&�d*�_0��Ʉv��h �]'u�o��̿{BGB�8����g����SH��K�A���9�҆��H�`BT���b��W�2�h���d8 c����`]�L����<��L�	�d��F����n�l����'q�6��0^0�8-�v���(��+,=�������w?[�8�˗[2$ ��ά9+��������j��`�D�n��S��J�i�RYD��r���fbE������yaM�Md^T|�R70^k4�4���n�g'���r�GV	�����s-@1�g�>V�����o�(iӖ(qS�e�3���«�;]*i�0휯v�K��3��_eCϲ�y�n=�HO�m5�C3v�HNA�&6�x˖�̄�`�f�$}�O��]��V"n���')��!gT���V�p��h���&����n�9�wy<_H�-{2�A*�0��h3���2��j�[�X�8<��	>�h�:A�"��_��u���R�o	/�Zp]�Jf8�
��`��t&fQ��RR�D�ö�Q2a�C�����t�u�?�	�򀑹}p{1����v�u-A/�oM��_�۟Y{u��P����^ҕ�e�(�DT#}�S0��3Ǌ��8L{�T�B��Z�T�䜂��`�5pRt��6Us2��l�>a� �-�Ap;����N�����i�yaנqY�P"������>[҃f�α�T���c ���9��}P�&��5h�L*�+���(�đ�� Q�j��T7�<"���K���jD�q�����
v��$W���m���8K�g����iHV�<����kũV�_A;2U��y'��LG#&���ҭ�����0`,�>�:rD�Wf_��e���Q��f^L8�Z׈\��1�q�{v�4)X@G-L!\5�7'9�.BN��G�G��w0�-��0��i�O=�5E5�k|ʔ�E�/��澥�$�SK,E��idjۃxKʓi�����sQ�E���_u��j��6�`z�t�Z����P��I�a���'��=����W6]��d��z���������v����nɫ5Jm"�*� _)���y_��`��30VQ�1VvzR�GK
����Oy�Ѻ��+c�d%>�	�1�������<�&�D�K%Ű���%�,b.�X�uks�-H�$����N4�0M���&���e)E��͐����\�X X=����=��~̓[�';|ޝ�ad���dP�]n�e6�� ro��) ���qU�W��#$BV�� m�5���zr����q�a(B��a���P����HP��<F�.�&$�=����)�n�8�Iiu��'@��~8B��H��ϵ���Ve��}ѹ�yh�-�'��*#��<����?W��������s�b)�נ��6Lҟ`Fљ�@'ɦ�'҆"����4rh?\�����Q"��-�߽��;�o_z$,�e��/�����i��@g�(8	��t���� h�SmUS��]Ȧ)H�8`$.b����yt�Ѕ�F6~'֣x������!H-R��J��y%�Y�#�k!O��R�=Q�	���P��e-�7�0�Pz}�%IOٷ���5��DH�I�Sd�N�GZ�Zj���z�n>��(Ur�F9�O��d5��k��M},92�NME�yd0�Q��Qb@��#��5޴F�>�Z���KU~���#���'��P�Ū
D�!@�eyM�J\T=�U���O�<�.R���cqs�܆P�)'�������D���|�$��瞴�������ol�~��;݂lrc�s��Ll[6N�WF���kj��k�pv��4Q����#�җ��gie��Jk`!):s���Bk�C���}w��R/�4{�:R>/�[���Ġ:�����_W��s�¢��ޖ���)t9�O��"�t>NC9:{�O+c'�'Y5�"�G#�9�g�"��!�(+��@�6�H���y!�]|�u�j��[�]�ݓw|DHB�X=|M�o�X�*�ɔn&o��	r�Tp�V۶3�4jU��A����A������d��Ir�e� Գ��ٌ��+m~F�}����m�٫�#����z{eoT���:�u��]�	S����]�x���