XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180<>y�_������5k�m���Y���4W��ڎ,���b�N�!�V�ʶ]�@$��K��-H��&�=��yE�,�15�_]/��Ǆ��~�_\���+������a��*J��"w��jV6ow+�	ed	�'��ntk�8�g����l��T�����IT���'�!�A!Yo�ܩS���7��JC��F�<��[�5�����O.ƙ�z*
K����e�8�@)���� �Agi���\�N[�I��"m�}�aU��ҕ�e3D&�~Fp�P�?�I��5���8��2ù���VQ�`1����S�� 3S��4��m�lk In-/�i�X�:��~���3�7�Kh�����R�U����.-�8X���a!C,��' /���u�\XlxV61EB     400     180��
�ގݙ5� �-d#^��*�_���y�Q[�Mf�1G�G�z,)<��ݵ�C��N|�j	����
���)�>��:��]�j�*����ޠ,�͐c��^m�L����է�וW�ò�� ����-�\��������c�y �V�p���l����џAf2DeY*\�������ix!�|�����8��.¯��r�?���j��Y�e�d�Z��!��K:��t��dӬ]��~���AM�SlWE���&�l��=�R��d��Iϣ[ۤD<��F%�:j�[��1y���� cQ�ö�����g'����{۸�� ����TH׀�c���Q���׸�T�~����,<ϭ}���(Ӿ�M��O~XlxV61EB     400      e0��}�eR.CfQ(�%QJ�$����6%}�Ia[n��5w`~FHq ��\���şAR�M�@ �6��p���x{U�:*�^���{�&��h���Y���
�x���c�.w����7ڌ��ce�''4��!��|,�{N�Ё\\ ���k�B��
�gb
k���:%���Au�-c���!�> �,�J�zbXEm�5톎,q������b����+:7F.���	XlxV61EB     400     140��K��3����s��0��`�l�`���Bמ=�����@�'U[8�<Y��"��O��U�&���kݷ�)<-���4t�)��ܠй:�7�_
���N�����в�LhUy}����V2:)�T�_C�#߲��� �7X��ꚸ*ƭ�h֦�u0>چ�Mن%��� ��[�J�Q�a&�ڙѨq8P���0��4|��:_/pS�c*����(�c��Z��-O�R��kA���@�Y:b!�X�U�J�-3>�+�u\���W�������*2rm�R��O沧���tU]����"(XlxV61EB     400     150�F�ٰwN�v���0�p�mw�����n�ɭ�ChSm:R씷,�׷�0;r��	q6y�Bf������}lr=!�-B��3�"��\���<u%K��ACC�J.ӒH�H��?�/�����i��1R�������� ���i��V-�m��(��_B3����؋��R�D`��H�����=���?ĳ�f]ϫ���2���hE�f)��4c�ܭχ2�tk�vw�18+(�|䙴�Lxe�尼�`)��F-��Zh�@�>�� �s_��ϝ�P�]tk�JR�W�I�g^�v�GJ���(͸Ԛ������2:߬�W���T�󌶇�@YXlxV61EB     400     140Q�����	$�.����s�����H�r׻���Lf��	[WhE���V��d��"]a[���q���h
m[�^���cp�5�G�cb�+���������qBZ"��rkiK�w�~�r���'-4����[4��z3Ib6�j�;�Զ��Z�,x3{�F R��V_���-Y`��h��B�n�5��J@$���8��Je��j�~8�ھ[*> V�C��0	�v��B�fZ����y�Í�9'���R$�����W�d��N��P�G��՗�d�����2 �hS'���E��+=Xv�k����.�2�'�S���~'��m��XlxV61EB     400     140[/

�F�`��Zp�U���~s��U%�:�?��~��lf�&���Bz&���]��LG8���J�h9a�v\n39.h�2)y�d��D�%�dC��1A���/���� �#R��8�#qViD��P�7�����D�r�zj#���#�4@S<;a���O��L ��?p�1c��������AD}�Z5rِ�=�Z�*0ġ�AF����~�Z:����m#��>N��H�I�Q��ž�v��p:9l3�)f"U��q1������{;dAp	�x�s~�$����Ñ���?@��dU.ih}P���l����O�XlxV61EB     400     120��aw������mx��fٲR}��X��R�;�M'���RR�Ɖ�����S�M��JG��`�Zo�KyL�Q���_��j�cv�i�U�[�HЛM߬�����ϴ{�|b{�f�A����t��>y0}Yʜ�` p�PG�5�ڤ�a�g��L�>�H%"P@�酊:,�)�|C<��@@��q�������J$�V�b����x��Q��Hr	����|��]��١�b�^�Z���QJ9�����FU�/�3V��aB��f��)�^�����3����p�3�2XlxV61EB     1fa      d0�4e�*����ݙ�k�^��r[�胈�3U�]t4Q�}��2��<��6��>tFۛ4O�l��9pC@�o��ι�8�SԬ�]�9�A���~�V��e��;��Og�˯n�$�|?�N���I>0�T�a2�֤)J���S�e�,b��q�6^���]��c���>D�}�.��v�2ԝ�V";�?fC�N�g,����U�