XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160��Xoj9��o�\����8d9�8���ڀA<��x�Êy��\����`2�'�D�� SxѨ�WT9kI��� ����Qa��d�0ꔓ�
z��/jr[�������+k�`f�o�]:�QՂIT��ZF�M����ᬹ��q��I����n\5��*�Rt�$��͗K�l�s������)XU�𷛕�v�]���o��ԝF��(t�X*`hw�]iLb��K�,X�C|��)��������a�e�La��N�6Ց���wF���q�]������4  �.HM�Y�%���N�A��Ù�Jx'Zg�?�P凎�~�n^1zy��r���AD�AG(3Ā��WM�XlxV61EB     400     100��/l��k���/=k�p��ﱆ��8�O���/	�L���p�V�m�ن�b�a��鼪'�ę1NQ{d�`te*���6w�J7��_�o�"�ZSHӯjI���MOJ�Q��q���I@IqZ�jL1[�3�l��@{d�+]�4p��N��+�^a�+����1[�!�^S-w�oх.~�ں��X_�QԮ���%�g/j��}� ���Q2�&���N���~��j 5e���Y~ճz��L�8�n���fXlxV61EB     400     100u s���F�zє���o�"�t�u��G�����)���>n��^�t �"�bd��~Χjܰs�?.�����n�G�иP�6�����+������_�\���z�t���b��=�w�;�믄U�Xdq������Y	�1��靈�y��s��+h3t�����.�`~�^N%�h�"�ы �qV	��I[k�55.�H)/�|(-:�>��/AL���}��{���<1�zTT:*hdn�D��|�P�s�/�.wXlxV61EB     400     160����]����9@e��1����M��t����+d:ٗ�:��c4�� :Ku���%�W0�b��zG)�*S�\�B�ίc=vhZ��vb�*2H���v�6Yq�f�:ݺL��Lӳ�虪��S!"��B��L�ޏV���ϖ{yП4m��iҺEA�b��2�	���H�'0-�D.HC��%	�(�X��'��q���WQN�X�	�h_�B΄��9��3���U��^�9��������Y����_��v�mF����ZeY�����A�ث�rlm���3�XH�^���a��n|ڊ9�;N��y�Rm�%3a�Ǿq�׷G��la~��=���wAEm��+��XlxV61EB     400     120��yy�V���}{Il�1�Fp![!���L��8�8�ލ��,S^�|q�B����
�~2C�9g#�f�~@�xȂ<��d_���� ��o�==�\��m4�Ѷ���J�]Y���o���0#z��W��P��D��Cy�$0Cn�X�<\�z�T�������K�2�L��}���h	&�:�+;�[&��;�k�v��zCK:����w�1W�@�n.�<Q�@�T=���X����%Ґs/�g��j�x�n������:;��m�.�����qc~�;�xG�HXlxV61EB     400     150��,���V �^�f.Ӎ��5���;,�ܪ� �u%��{��I����B��$]���o-.��Q�����DM�\�3�.m����YJ9���4� yH��[�2_�*?����3{�q{�#�ش�%���j߽�}a��b��C���,7���u����!�O����F�5X�{(��=(3�d�т����<bO���D�W�p�j�\Ĺ�/�F�ZѪ�D�no3�s�! �s��2.��h_>"���x�����+>~|_ڬ��/h���hG~hp�o�ij�@�th�ٷM�3;6I�:p_G�� X!':���Ns�2��X�|�'�n�NSH 4��XlxV61EB     400     110�i�} ҽ��8VQ�5tNd�~.���g�}�?� �OGܰ�����)��Ԣ�>��Y�jdNe�܇:ڵ��Ed��5�����l�=Q��TVY��IUTH��L�Ue<�K��1'y��'0��ᎆnÅY11�6�EW{�~�قR�#��-B�9j�o��6K/��W[�E/�[�֕�>����n�e�7�K���@���K�Q���d����=�t�d0 +N+d�r=��cn��+!�N��բ��o׶���toԩ߈ .�i����}���XlxV61EB     400     100�b�:��-�Τ����K�c�9/FH��?�sƃPD'��%uc�)�]��<��XKX�tc�-���}�ϕ��2��J�<��0>iU�NK�?�R��R:��qVB�c����Ub��_J<,Q�cc�^&�9@����z_냵>����f��ȫ��5�O������ Y(�Ojǀ�P�>��_���ߩ�bj�zkF�����KK0�6P�qd�|.ީ�f�˨N���N�gD����/�iTbb�A֛�i'M�i��lrt�XlxV61EB     400     150�)&x.0��HPf���g�p��%b���QwD�ƶKd�@�E�7W�M:t��p�1UK�v�P0�s�WHws�'����8*m䜰�����\�N�_\�	 �G�x ^-��i���$��FTRz�"���%*ŖvJl;���!��ح����*E�̰Y"
�>�K��.���-y�D��o��/��v�OC��j���ެc�g|ƁWs��b��嫞���:�[���xn�zԽ�3����K�(#f�u9�mfxp�j�lC2��|���P%�G�V
LSDR@�X��	�KZ��q.��\�,�� �ܝ�{�AYahS������7�7)�@�\SXlxV61EB     400     150tSo!��?��{F�~��I��uK�̪J�g�0:��h؊�I��L�;�cx#��ݰ��s|,b��i�N�a�o�m�М���4K�Wi��1DIϊ����	zA!�2��V�L�۩ぱS8�=��ihlV���l����!��v��B��*j��*yB�������WKdO=�S�c�+�y��J����&��z������r�$v��Շ�������2����F
}���:c�x�#�����*���tj0&�E�^48��X_b��=9T��d(�.S[}�ʙ%U����%l�kO��m�J�mW�S��2���GG�R���g�XlxV61EB     400     140��$��B���0�"�[�	�U�q��lsN:Y���oF�ZKN"��i�&��"��!2�BF���ͽ�S�S ݷ�{7�T�R�X&.���s���Q�4���~�"�BN��GZq�ץ� 3�	Of�C��j�_D\�F�q��D���"��Ǣ�y.��Qm�������0ˎ.�Q�\ZYo�IdI����<"�ds��E��18Xq�ˁ�O:����5��GDm��$��$,8*�BS�%��-0aS:�E1zId��^������On]+6�(�Z@}s��-�9�<�~�y��f��UD�Ь���V���T�XlxV61EB     400     190&63��Q��{&�ǃʟ��"?�[� ��jQ�r-��\{)��Q�R�C2�g4�%�lxo �̝�t��x�J�@c��9%�!�k%�\�c��|(I� �v3�.��砣M{3����M?%Mj� q��
ú�FĲ\l���αƶ��2^j�_~q��ſщxݲ2p��sJ�8�sp����J�'����Z7��î�f{^^��s�Z|���1۽���k^������=����g�cG��l�b�_��L�AN��P���g:��;A����T���v嬻��𤋈�d����)��N���Z��V�VK��ڎ^�:�Tn��V��*�l�-%I�%M�JΒϛ�yx��f�3���ȏ[!���a�7j/��T� �)����Ր�RT�h��XlxV61EB      81      60C�+��0e�����*�=�A?���!����z&e+���P#ȡk<���ɄmT<�s�I0&$ƀq�ڂ�d'�y�G��0��'��*��B�B^`~�%