XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170rG���8ܱP�ݤ�G3�~�X���-�)���Ix���`��<��S'D���k���ʖ�if��0�X�FG���B�:�^)���OF�j�s��	�= �����YK��uM� �dqe��Us��-��M�ޓz���i��o-�A0�_���4���<C�T�C�?#��j���5���=�~�1�:�R�1�Q�-:O�ޛ��ù�v�ly��3�P���7��d6$W�*�Y�Xp��G��\���~���'Pj���_����+&h�{�x���x~%�_�.�05�'I�R^qK�jd�o��@ȗ��B��K�Bu��TQ��/�=gI�+��������L1�5�6H�Դ���#��h�PZ�f?�XlxV61EB     400     160�Y�q�s��P��U�����,�4�rζD���4�"d��B}��3��>DI���̘-��.ZT�S��o��A}���2�|�K�����TqC�^q�����od�6�b얷1W� ��(�}mc��Z*���V�dϥ]�T����j�+z����'�-��ƚ�E ��SK�u{8MԽk*�l��p'b\�?t$�2C!Zmͬ{Y�h��S:N�͊>\2�,7X�Άv��b?�����4��T{�珁߳$pB&/��H!ư�~i�Z��\ݲ���Yy�����ӆ�������p�`Xٛ<��"��(:3�[�b7͹sx��'+R���#���?o�'*�c�4:��XlxV61EB     400     170��s��t�ĉtԑ�U ���^	�� a`��Ir#�(�#����`�_��=�<���Ye���7������9�D�Wl	#�҉D�o����2i&H8W߽ﺕy��5 @�۲K��kz�>����-����>��d���1���t���GF.�Vs]�9�o���ݴl*f	��v�v� ���\#Q|3����b�u�F�i�K�𐱔l��J��\T�q�~�E�!$�bN�,��n/��?%���@���:F�D�[v<ϻPQ�T�r�g��H;�P�L�ĖӚ9��L# ,������S����R�le��Гjw�[�Y(����E�u���:���
A�;��xN��pb�OT�v����NXlxV61EB     400     120����=����?l]�ݔ/�j6>a)��}���%m`+.�yGSpb!�{d�� �����Ma�cL���)o� ���f�pɆ4r�?ͤ�Ҋ��cW��aU�I^)��@��'���TǾ�K��/�#^���4e�H�#�_j)6sںDv8�a�ǻ�lw���4���Ӹ�VdLM�!�kKY��i���nJ���DVr�-�/�e��e��n�n�`�9FT=S��YM�0ݙ2��#�!�Syﳰ�HR��l�A	H2����TG�_�+^��=�1���?}B�+�pOb/v@�XlxV61EB     400     150��یo��$S�[%����܆��y���C<�r��Z"��⟗�߆�w�e���XO9=�T����ѡ���dnh�w,Z�)|~���Aژ/�.^����F`I��#1�L�Ƕ�]tg�P��ి�)3o��b��@���� =7���D�{"��6��rՖ&i�\�G��V�gw���I��I̗ۮ��
�!�b*W���r$�.�e�ќ-4���C}��~���r6�H}U�Z���H�y�Xk�cl�r5]C�|��(Hh���
�p7�������_+4iBQ�g�AɓnO`.�R���X�"�<�����_�wN�Pr;�#�7�dG�`e?XlxV61EB     400     170�����p�1E��;�qs*��H�՞�˜�)�����qS=�s]|�{��O���(T�U�,�k��ы��~�Hk��X"���Ǟ�MƻK���M����#��{���$�k���R�*h��m�g�D�A�Ꮼ��hg �c�L�	q������0��3��Zg��K��P�ܳI�=��ҩ˺���S�T=�W}�2{����p�O�{�X{��(h�?"y��t���[T�Õyqx�K��r�Qr���l��/�+h�u��^q�7U݃}�a�ē�hMH.��&-��n�}A2��!�/Q�p����۫o�P����p�e��4Pd1z��e��-`�����{%�;Ru����XlxV61EB     400     140�}��#S83���۳;o��AĊ��<JW����[6W��Ǫk|/�����ؾc��$��a�2��\Vq2��jc�~_D&��<`�x���?h��¢������u5i��{�>�S�Gݒj��
�����aq��X�j��#o�
-�H2qrO喝*�K"���OW��k݋>e�f�!��q��Q�nٹk���˧��E(�.�8Sp�<�y��[�I;�4�2DT��3�{��E'�[%�����.��0&ٱ����*�Ύ ��'.z���uo���Faڃ��G\��c��1�fxN14ֺ�H�2��E9Q��XlxV61EB     400     1b0s�]h��cÄ�~�����Շ<�'�&�AG-�!d,�/�WǧF���#�W[���G����Xg�yPu��+��/�q/ºw'͜d,������U�I��`� ������VTp#-�KC�l!�e�C>�l@�7̚����j�`.+A#U݅K��eb��B䣁>B<Wh��Z� X��>>n^X�7�o���4���Y��<�x7�GĹsw��`��DJ��-�O�J
�)�D��|'�_�W�n+��LI*���~��`�)S3OV��x���X0���x�qg`i�����D�iN����]�O��ng)sYqn� Ci�i�t� /w�eu�;��@ݜ�M���2�M�L~�@�X��r&dw�����^�������sL�H~ܾI���.�4�Y0ڱ�em�~�|���:;��ɥ�m'��>� ZXlxV61EB     224      f0�W�r@}��es<�$|������6>|�q�LĒ(_��,(H�w�D;"��X�^~m�j�8ˤ��,Y��<QZ`��iɤ�<���цr�<o羊H�"���H_�{�|欈��͠)��ҵ��4�1;� &j ԤT�m*�uݿ����Z
�p�dP�A /��6�2e54��]>���M� ��ߜ֗�Ck�]�`{��M�l��^7#������$��QBH3