XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u�yf��)n�x���l�x �5�-%��_9�s;*��k�B��ʥ/)��A���Lf��&��(�,�p��?�q}d��y��Xx#��5RN�ʳ!�_@�v8TyWS#*޹�懒=U��]IN�65�V���p&�Ɲ�2,��,��5`��w\~B_pC��S#����W��`�q�g�G$,��h�y���������y[O��}�����k�`jb�Ď��F� ����s�Y��&?�|Mﻕx��+�@�zX���X� :�zn�;@1��'JMZ����ɵ!9�aP������m��iG����#8)'���vo,�Н����(41��AM�v��bzo�j٨NP�a�O���x��ƶ�_�����&�ۈ���o���!�P��P�B5K�ZT>���I@�=���$�m+_�S��˴B�A���Ѹ�bH�BR/���b�}5Ұ�_��N����ޒ�H��n��gH�_3s�w�p�&'�C ش���5���}æ&�f���A���j��DX�a=�}�G�H��-C��_��JG�ӑ��4����!Ǻ�iҜhR�/ �Wv9{�L��W7K��(������.X�O� �����|}g�3�$��߯��f��K�`q�Zd!LD�E�@�3�1�q�h��g�O�j�Хߤ�u/[I��X!9(B:L=����_��B9�G�~JŁ��	���ďl��2���@lk��& >��m�[���Uߛ��cd�_��e�6��A�����QvKXlxVHYEB     400     170�w �j�2�2��h�0*�+cN���G�/o���U�]e�l�m޸	jD��$�*Hi��'Ɋ�ߠ(��b��3�����F�m@�������sޝ�(, �����	$�\;�,#Vz��q ��R�홺�iN�IZ-r��[�f���D`\�!�=:�Ӽ��k�WNŀ~ �Q�#�,�~�UQ�B�YIV�-�꒞���/x�}@N�j4�@���:��^w`����-��R.&{N2���>�
�/��%�j����-�X��o�	����Xym�P���0BYѐ��q����������D@V?n��c�P>:3J��d���66���(��S^�<0�V�բ&U�&/�X� `?��+��bk�XlxVHYEB     400     1b0>�Ω�ӻ���NJ�?s�i�4��w.E��]Z�]Ohcy�-��M_�>��r�M��m_�B׍ґ._x���V�2���]��8�u��)�8և�
s��Ìx9��̊[8��S�ʗr�UR�h�9�%CLv��@�m����K�a�i���-q��=:s�'L�Et*�U�>�)�o)��x8@���8�gQ����E���X�#�
����ڠP��q���`�f"��7��D]Fv��	9�g�C��15�)�I�F�=�����iy�чN� �� -�h��Wy�'�{�����ą��@>�O�I{4�S}�Z�*�OR2�%x��n���K'��f�~;c-�G7�����+�+��:��Ds��7��o�!)f��g.�b#����)9.>n@�k��)��X sὍ2c����5�H��o�u�&��XlxVHYEB     400     170���侻��J3���*Z��'U<�@�5S��$J@��͠ (1d��tcI��X��� ��m7:#4�P�zIO��\��<��B<$��J7k1���b��p8,Y=�,n���\�o���|/e�"����`v7=6��id��������!���)�}H��	�uϋ����t��g��׭�:l<CHR1h6R��*��gަ�Mh�C��k��L}�� �Wal��~�`0=d�rzr�.�$�J���#�,���VՕ�Wt�)3�ߞ4���Y�c^`�o���V'�<DU^�=`ߧ1�_�gJ#=TW�^o�&���d��R4�]:>�� >���6���a>ҍ�/z,<?WOx_5fXlxVHYEB     400     180$��NW5�!İo9d��df�a�"/=ˮ¸�0籎�D�r������%���4�&\%�dA�LX�HXg�4�Wݾ�� �f���g-�-Kq2�=@$��_H)�Dm��-�}5�'q��8�A���I.,~�Y�v�p;Z��RP�$yOǬ�� ��2�{��E�kJ!�!ӿZ�C��x��媼��1v5��. ss�+I���
˿�r�f��ꡁ�N������&*}����˿��v>=n䈎��v�J�����`���S>�cy~xc�*�%�v+w�'BN)e�zr�����\e@���w��3�P7�� @�6Xo��Õ����vs"jv��zE�=���t����8W�!R�1 ���ʪ����}$dV��瓼t��XlxVHYEB     400     170!����db��Ol��y��XB�ÿhA�>�m*R�z:Z�I�Z��k��Jo zc=Ͻ�8c>E��6�7�#��o��������`ż�gn�b��^� �i"����������2�Tr� .�TmN
��JƎ��u�I����8h��Y5	�o#���ɇo%t�����鵻�S���6n�E%�x��Q��IO�r5҇�o�7�A����z˴.4�ٛ:{Sr����g2oxH-C�D������Y��k5��))߇��@�}j��D��B"��e���1Y� �/Nh�Z�-HXB�7�7-�ŀ����7n�	�Fu]SF�B�!�St~�՜�����I�����,�3�� ����d��#L2 rXlxVHYEB     400      e0&,��q["{tq)���@bR1Η���'2���<��Z)�Q�T�R��lU6_F�F���H�v�z#C,n�X�;�j���5OT�
���<5єe�?+��o�V��N����s�__�����[	1ED�)<���~�-%��NҸ�O�T�y���C���/r���4�w- �X���O���!V��P#0
����QPB"�űr�=��꧟���wJ�XlxVHYEB     400     140Х�"����,�S��U),:�(W���������6�P�̪�|�$٥�}B�L�q�R�.������)D�wV�!�T���#Wؤ4�K�!��ո�b%ޜ���c�6o�Y3Y��o�kW�T_�EIctԸ��=��o	I�[ l���#˯���&�!�&����'�*s�O��ʰN�[]>)��A�-/%*-���}@�L�)
"�#��J�U"?���|�E�6�&�E6�:�f�q�V(�(;$�tG��̖���v�I���IX��(���.�P(7��f�v��ݺ
>a2b]����<Q�!�>�5�cQ�V�m�~v�n�XlxVHYEB     400     150d��jCj����/�`�υ������� ~�8Iˬ �67QX���5�BQk+V7�i�S|t�t�[��،�C�l�?ސ����< �^��OɌs��g�n�l!{��)�7��31�H�;.���D��\9�s@�v%.B��'/y�e��~�����vC�2����VX��b�P�Ց�Cs�J�@���a�޾G�+�w6i
n�t����+��<Md)K�}҉�GL|x��������n�9G+.`�[Y��И�|�kw��|sb��Io��\|J(���N��`��;�/ub/���]~V_������u�h�*���m��06�XW�g���o��a��`vXlxVHYEB     400     1800�U��H��B�;_ļ�ըs�|��W:��0x��*��������5?B����}$��빜���#��i��觭�s�> �l��I���%�YX�n�7(��Ѝ	5�I��%���c�'� �<�=��2g�1�t֖�Kn����c-������J�߇�d��A}��H�/��͸(tr:̷~���vXs�x~�a8Vh�=����>��C��|XC�mn��
����()����{^�6ӭg|�iL2[�S|�mf�G�  �
"��W�%����PW�!*��1S�+ ;(�H�P�'b�x�{2etۓCN^y��i�6��X�)�H�!�u=��e-$����'������O�5�a�_=�C�XlxVHYEB     400     180����Y/���H�H�Q�7C�p���啧�H<oH����$跓q,��D�gO��Q"'��~�y�4-�,?�!��ω��D���|.	.�aX��s�E����f�������^ǰ�p�>q���(A�4�"������sk�%#��}?6�S4����7�e�\�"����L�~�Pl �SAw31��L����z�|��W���E!���b���"'��`�A�T�jTE�);�`����c��8��ITf:�>w<,"��#�i�la�9����؉L��I�t� |������5�u+��p�� �4�}���.�GZ�\�h�Jٖx{�}5�}���_"B�/�-O���S������ƭ�[�XlxVHYEB     400      e0F���|� �3xG�[CjF�!�-�v�[L�W���sYج ��e��x�"��J��w�~�y�D����V�_ў���J��Ɛ�U�,k钓<�c16�/)Lj��>��q<s�k��r�ӥJ�9?4ܨ�՚��&W�$��$�s���V:���0�q�E��N~�����Z|(�؅cv\Ra+^L�Rg��,�jЅ������osx�Y���EXlxVHYEB     400      b0{�w��3-ϿL�ok��k��������)#y����Qc��S��V'��^i&fx�2h]�n�w$}<_��Y��ٵ�hhcF����Fbc���NN0K�8��"J�A�+��q���{��������.a�=��6)[��]�F��J��/�g_ג��P_������VXlxVHYEB     400      f0�ȧ�)�rHL���\S�D�>Wa�N~��Y��fM�%�千A���团���Xa�}��Et�d��ל��lV�6OOn��"�/;u�������v�S�yr ��b��AN����Ь+�\8���Qb��*�{�m����^�_���_v�#�Ӻ���cL�8�� #DC�S~��\��#:��eʶ����^���'����1�2i�ǯ%~d��Ɠ�6�w�2��HR��+�0�Wd��XlxVHYEB     400      e0P ��`V˔}�C�h����rF��
��T�e����N!�M��X�1.k��͉�	���b||N�����*D��-N"�u���#j0��:�Ed�ar��~^c$���*!s�Zea�70�7e��κ굣opJ`�9�<��|���C��mr��cAf���h��{�����埽Q����V٫f��^J����,q)�l09F�':K�9��0�XlxVHYEB     400     170\�%^^V�ko���'//b��5 �a��%�O�C%�Y��B��&q��^wzݨ���]9�r<�%��|l�r��T;�Y�������3�c��%-%´[Y܄�I��!� �m.^���N�1m��`J��C�.Y
�g_�Aw
���.�x�P[?fK��ɛ*�-�4��)!4�/�Z�0��Ƴ$]]�C)�9�*�JK��;�Sv�ʳ=("�\#_�(TOi�t���=����ҭL?�	�-� n�5:�u+�f�s��#�J�&�rAI�D_V�KX��<@��CᨖB2Z��:e�gNQ,�c�'�jYv�ˆwc�L4ۂ1{�-�l�C��-�J8d�	Hh#�eI��d�O�o���>����XlxVHYEB     400     130ܰCNf�%c�^��Ӎ(9P�76�/o`H~����׮��+�ծ�(<���ur.A��"�R�.�b�>?�8-T�P����s;�"���}J�ٔOg8g���̆`�m��� �3�;��9a��	얛>D����W"��SCz�LE������]fAn��J���F@p������`Z��E�ȱ�"c��}��d��fd�ǙYO���a�Nɱ�`�7^ʺ�n�v`;���Sr�{c�)�a���1m_WQBˬ�ґ縸$�G-\P�����e���InuNU<;���O�����?:9|XlxVHYEB     400     110P�Y�v�Oh	.SyO���f����R݌���CD�]ӂT����̃%��y� �
�E7�F3�dGqՎ�Z�q�4�NQ����u@I������88K�^[�r�Jl^Ȃ9?o+A,ƨ��Y�!6�5�Kz����[�����Yw
��Lcj����4�����W�m2$�GaB|�	�=�QM!T�|���b4%mM|4+�,=�i��'iL?'����Z�2�Tn䢤Y�4#Z&�ˑ/dg�CB��akV,��q�[<�ѡ�b�����Ε�GƐXlxVHYEB     400     150M�v���'9��}����5n�m���&� �b]���3$��pu�z������-���0?�1�4:�O_[/��嘇>�/��"VV�Հ]�S��2lK	�Ip��d�y�Gx)߁�wsf�pC��@��>1�s*�IA&]@������e�C��U��x^l����&�{�ydo�bs����N�SZ��H�Lr~���@�����5��
�>	��Vn�Kv��19�y����	EIŅ�=��Z:��������p�,��vƨS��������/L�p$������&�Y�����jIn 7e��E����TU��j%)�(��M�^�� ֠+tXlxVHYEB     400      b0�'�����^A5ٚ��+*%� ��X��c��� t%2�j
�;�ϵ1}�T��x��K,L'�avv�����2-sZ_]e4�`��\���9�z3{� 0:��O��jU���/�MU�=n� 木���l] !�gw9�
��"����=ǂr����QCM$"� !��XlxVHYEB     400      c0��l��T�B��yL#���)J�UDx�\�SA�HO*����(y��87��4��[@S檦?<�VI���R�8P�|o��؟��brʺ�.e&��Z,z6soI��� �U�f�R��P�wY�MK����՝����-��m�L}�\�n��h;��s*�SD}�ㄲ�?�6��!0SUK~���XlxVHYEB     400     170�oK�،�Z���5#	j���|���ٚ���h� -�:>MF#�bз�V;����-��)�?�$��ml=@n�a����Q��bw�Yx�@hIv�#[`�DɈ
�֑�5���b4/��I��L���BC���\�����B�C\��H����w������&�a���0հ^:�����1B����7�ٔ���'�Z����<�vy��_�{�N�Ox#V��]��۞ݘ�g�_D�َ�	x�6��&�E*�u�U^
�F�DrQ�c{�V~-~w��f�k�_��4C)ntK@W��fw :.�S�]���.F�]P*<~F3��ú?�o>�?P�`��$ XlxVHYEB     400     190���EZ�n�h�z}Ɩe+�� �d�L�`[$]�s-3����T�Ӣi��j]�/'��vk&�L6���Uu��(br?,@�u͕^(~������8��F��" ��9:6W�@���/�{�%��b�� [�_�,�����f)�-;�g�Qj;��)Φ�ii�뀧ҭi��*�(�X��ě�c�Wǎk�|ɪn.gu����� PO�f5��D�F��u��� �dɣ�
[�7V��Jh}꘴l t۞�����r�Ǌ}�5�1��ʸ�p�����h7{�g����	�pl�}ǈ�����=�,��S58�	���K2C�h��n;�>�:t4���QefR�@��b2�Z=K?sco�����#�?�K�����0�b5YHr�g����p;�XlxVHYEB     400      f0����:�<r~!�)�mc{��z�S��&�/�L��ȝ�]�]���D��qK�u�G4�Ȼ����6��c�����?P3�躕�J鑓"=���
=e���_:OXm!��;@�.��_���O����c��]:�U,E�׬æ�D�5��C{�alM��a~ F�ܝ�<_Z����a�l9`|����Nh`Iɚd�O��ʞ�|_c�G��w����A������{�aV�Y�XlxVHYEB     400     140�S���0��_Ȉ\��M��<vx����4��N�t]ˍ����ޅ4d�o�!6�"�ZMoJ[��[[r�a���:!���p�7e`�~H3ߐq�/�
�2��>��'��wm���7��9Yނ->���m���L:F�=.ڸ��^b,k/>��Wt�� ��uP���!6��DnI��-8�/G�b�� �}USA�a���C�"�,��2���OP܁N~Z��em�Һ��8(�<�d]�σPX�GF��D�����Gh�n�
��-�y�jmd�U�Ҥ�s����vTV'����O�m��M70(�XlxVHYEB     400     110>��;h^t����겎�z$Š���2ls�4�8T���(�\ױfW�a8��~���A�"I�� Ht�5{��r�L��|2���K�wM��,��Yt("����Ō.���<�����;'�~ 唶y�#F�������#���>�JP��� ��1r3Z���n���1�x�9��������,��Ô�T@�����'	9��,;:R䭿P<#%�f
��y�@W�M�q����:>���H�:�i�ػk��5��� -ʞ��18�XlxVHYEB     400     100[r��Nr�uJt�S�ʎ��Ŧ�	�aL���#Hq�F��U�׌Euߖ�#4�W�Uq$�mzX&�O"7�#��=�we*���ȳ�%��Kza�m��!�#��8���
���"m�� M3�	�F�O!��ӂh�qtR�gc�I�ݬg�F��2�y�6�q�s^{v�6\�cL7ۜ�lh__@а��6A�Ӣ�>�������4<.`1�$�������*پ W��У�s��;�D��_[j�l�XlxVHYEB     400     110�6x���~�)���M8�3{L���p�o��F�<�tma�fV�Q웞���J= ����#��d��	��\%�,'R�<Evߩ��d�������ȏpA�P?�⬚��Q�`���(cN{�HT1V��\0��=��]7�w�C9�
��Uz"�MA��X\�F��};kͶ̤��T!�X�,��H`,��D_v9�V�����|gZ �P]o��\�N�acNE-�Ca�c�Ť�J�%d/80��~��\E��U){�gjȕFXlxVHYEB     400     100h���6�v�8 	s�T��fB�;P�8�g̹	WN���qDىR�V�Bt#\����Ss��"@�Q�VFA��q���i��-��Cʢ���m���܅2	�ͥ��|o9D`w��Cf�,�*h��Md�+�R�G.Q/i���ȴ!7q�G 1l���	���7�z��f��*)�s��_�����C��x�3��������H?F)&L,�L,�u��0>_X�1�v�� ��CW��D~PJ�mQ�XlxVHYEB     400      f0?�eMN�/�0�9R_�y�w�Vn��+�L�;�|D�m�$In�bޠ��<N�Zo[���`��I�R9��8]'���W��<��x�0�N^������v?�h�䟌��\%"��)�N��
=7�`;v����x>o[���K�7�q�Y�t��� �'��,��`j�&��H|t�����0�~��ʫ<)wYgo��&qFIed�4A�u�s��Z^�Bd3Zo�Z+�Y�^ /��O��;q;���{f�XlxVHYEB     400     130�Q����u�]� G�$��b��W��r�����Q��Rj����:]E� �a���6jN��q�8m��.ߌB����Q��ˆ�ڪ��W4i�)�*�ut�~��e��&��
�o�_�x�R�x��[�*���@��B�0�#�6���I�}nX���}��1\B��X&ڛL��>�}�\��J%�~8ϵq�b�9��j���fz�3�-�LL�������t�3 5ן[z�C 3k�4�t�j�Kr�S��?e���y�O�O2JiYE�!��<�42}nJO���x/È�,>"�i��ҪXlxVHYEB     400     1a0�C����C2�1Ҭ}Ne��!~la��=l�O�/�k��[^H��[Dg	O�y�MG�]��Æ�z�;q�<�����S���G�y��k�%�c�FÀڭ}�4��R;)�Z�	%��YrۆKou]x�.��5MY��fQ6F�5S�S��;�,5pTqW�L~Z���G(���*-�JdF\����ZVl��M��>��ST�NO�P�F���`�6Q�r>���g �/�z��j)y3l%Ҟu7��r,Jz3���H/T�v��f�
O��Ƶa�	�Ǚǉ�: p�^q"��P5{{�\��
1��t�-��P��.:� Ǡ��v�'�*�wyC�������������h�Ie�ns�W�*Κ�����[Ω�����}��3ɪ3�m��Ľ`HO�����KY�FyXlxVHYEB     400     1a0u[d�5� �#����N�[7��_���M/x�O�l���������雼��U���
�O6��1�[ �4�H$Z�<�z4��6Źs� ��C�V SdáIX���v]�%Ɵ�#Y.����ԩ�����t�Z'-��#qp�0-�7����s#��5�\�u�u�
���X�;//U+M�jd���~��`�H��f%*�k�d��f�\Awz��k^P�P��^Md	E�;��&��S���᪱T�V���q:bv���ʰPa��Y��Q��f~ �6p�e7}]dx�������
H2��;Ku|ޙáhkAL=h��̠�l_G�(ٴ"C;�w�82�(��b��b����Xc�<�Iv�w1���k�R���jde�=j�$`���T�, S�#7o0_�'|k�Z	�7��XlxVHYEB     400     130:0e�\�AY�`�'�>AU�b��u���Ɠ��Cnr�l��T��21cy��Y��������.�=6��G�8p��9�8�1f�H��8�;�G>���UŃ���[��"�u[Ĳ�d"7|L n#��w��ݐ5��=���h+���h_C~�Ęٞ|�Y�+��ˤ�ڈ�C�pCG���S*�*��3W�6����jLƭ���ڪ�v�B�:��[���1L�U���3M%Nn�dxN��魞,&8q�������ϐ�$�"��Z����~��#bc����S��`���C�H��4�)��XlxVHYEB     400     150Q���8a���oj����a��
V���e�
�wV*R���;
;�Q�6#빙���&�}EODP���λ��^��U���S��^)��}( d	���2�Dဇ>�2RU����;�SVd�&�^��8�ma�TE�Jb��	�@g�D�~b+L?6���L$�7?���<�8i��hG_�g85�9q����>*�?a�wAٰv�[�j�	ۏ\���pR1�	�Z��Š��-i-���^�]e(ܽo���(����׭Oj$9���:YiUo�j�\��xY�?P�E&�Q)RܱB�d�����o~��b��]�����r���8g1XlxVHYEB     400     130ջ�DXf�"�S��]�$ՒB4��W��h2�;_P�3�
C_��z�0�w�&����g|��2��F���˻&������84�R�|p�����J�/�Z��
8i��+N|��9�_���ʦ�
sz {�>�tɥ����Ѝ��s7�8�R:��7���V�L�;x������q��P�е�.��h	���#��p��0���9�B<w�T	�n�K]VWW���w�[�a�<�q�Q폔^g�o���A�K����_~����[�� ���m.�6M���}0 �]�.F;{��5�guXlxVHYEB     400     160(G�٘y�ݐ�	6��ST6�eE�]Cۏ���jb2�[�R�-���uvN�N\����I/��WceUT�Q+3�c~U�D޴`\oW�Xo�(��_PP+gz^ s_��qmS��I��T��-⷏#��f�oEy��@�gq��/(ӂQ@N�ҝ�Ǒ��$�Jq�k�J]�z'd}@����{��*�:���W��R?`��-�×[���1r��ےB�o���$�헞"ң[�X�2�"33FE�+"OMۀ
GyՃ�n{�1����}m�2<�EXI-����q=���>
P�k��Bi��������/��I;j޺�C8��+Ie!��B�M�o�|�c'��	XlxVHYEB     400     160��f��S�p����ͮ[ۼ?���`ɴ��)>��ә:����63{��@ E�� h�'C�l�^<}�2�Z��R���V�7�&��V�`頇o��-漶Z(;MZ���SE���%(GU�f�7�(�\"dc�ёV2nX2�ox8�B���J�:?M0`��Gy��j
>ȫ���䠌�.u,��$��eJ����k�33O�����ܕ�;7���	�T�+�A.=ܜ�������a`_Bs�?[���v�x��B{Z�i�NO��Ld��
���7q~bInZ��s��o7����_�	Ѳ�O��N`iWb�v0l�ݭl���'�.��|�-�ʙ�u�0�a�
z'U�2(M�<;~�6�XlxVHYEB     400     180+]��B{+Be�;���i�_���"��G�˄xU���������v��L��ˉ���!�$��	r�r6�&0h�'�e�Y�-maAm��j�aOl?�G���7'�qIEBZ�BC�*�3.��^���֎K�"z	��K�a�2;�b?9��C��̏�֧����&��n�e`pV�۽j�0 �x֮��a[�H�*��YD��>�RBW\��
XG8�O͎	!/u��LxҴCGg�<�aBP���P��$�҈��ⲕp��&�WZU=����O��)Y��9j��9E�dL��Y�x��*Ji"(/;U��X�(�by��wdU6��yɔd�jB+�:��,��<i&��v�":�gT�����&����A�,�f8J��o�5XlxVHYEB     400     170
���>/�łV�ǻ�3��֊)�r!�}�����ۮ�L�]���[�"���u��9o�~���nf�K�>�"{uʴI�t4�?�.;�@5;�<�!k��4�#NM(�[}���J�i�����Y��OW�E�@
V ź3����TbF�&f�B�pF𣡈�Q��e���ґj�.��N�m�6��(G5 ����~.��93z�:�+�G4lx��[w���(̶�.3��'��+I��	9��6	ѱd?T�-���R���r�9�]��L�0^�j�f�h��]�V�|�kR��<Ut�������_����}��fA,��X����֦%zM���Z�� �ɄO�'4��.�8��:�������(��XlxVHYEB      7e      60Er�V~s�cA0��x��s��G�~J����nuY6�6���1N�^E �oEЃ� Uh$Uh�d����5_I��M����g$�t���Tiz��r