XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     150u�4G���h �;��H�NY�0� e�q0�fV{���A>�� j~���*X*zЦT�I�=�%5����g�vv�p��4���?�"�w(��.���`�]�<o��U����{'\p_XK�i;[�h�F�;�;!�А��ԧ�ApjLWG�	R�j��n%�^�.�g/*�CgT�b�K�b���{:�!�̸�Qr
�o�bpف��K7>�`w�ن$��A˭-�G0JE���]K��፱�L�Ѥ8.jK��|d ,*R�o��g,��Ԇ�[�P'A��_�Č�<!.d�B�jhbx4��8����J)�;����C����a�4��զDXlxV61EB     400     150[���a�.��9����?�Dg�N?lnA2`�	�:Y7M{�!�(cELS!.Xri?W�������79�	�(���VNGh͒�~�5����oX��!�9� ؛��ˠ��
�u�l������,��	�g���U=I���q��?�$_�Jb?r��w��c��]�A�S�~���V��9�;�N�)� �駄�Nln�p������m7�&VWد.���Ka%�J&�&�:I6f�uxU���Yω��A����sV��xx`R5j\,*�;�x4�������K�`L�]��U��i���~}P6���Uh�U7�呭�7|�ܔ9k>�XlxV61EB     400     180s��z��?�H�&��+4vN�߮0V�7�o�E��#�tene���Ά�[%�^���S*�2ݰ�xb%�v��C��p?���zi<�W�G�\�bQ�GZޝ���\�K:���t zG'�f��v)�\`)(�ޡ�y#�X��G=c��ΈT(f�d�����F3w#z�)�$��j2�P,�� `�l�&�~�7�������~VګV� תcĚ�$kڗ�z)5S�ge�5'����`��f�:�p��:�&�[YKP��/|�7�����DՕ��
#Q8?����ƻ4HKv�XlIhơj6�����_3�]��+G��L�z�LF�-:��>�ER�Sur������t'���ڲ�C���n�q��_?XlxV61EB     400     140�~*}R�)t�H���#
�[��O�U�dޕ;�-ң֭��(����
�Xk��Sޖ�O�O��(������J�F}	�}����bXt����V^�L|�K���z���&@���[�X�nhۮ|��v]�n4kG���7��^��!!U�/C*O���w�Rr���H#@�?��aCհ_N�1	�����z��k�Q��\�s��/���p������;�TĠ�.�w
)�BS�B`�0�w29�q �C�fA�x&��X��z�dQ2^"o��ȃ̖��ӵ@�)�K���Xm���wH�R��ˀ��]XlxV61EB     1ea      f0��Y�S��~0E�	���m1�R�8��o9��o�¢�t�B��7-
�>��V�%#��#�_�9<�,cH�_�GF���vȁ$	�y ��S�2*�.Z��'�ڿ��o�ݩy�y��,�Q$Ȋ�'퐇@F��!�>�.h֊sL�K�@~^��}��R
;8r׽H���s�����'�ƷM�[	��U�ګ릖�H���"����j�έC@���ڥ"�6�}����R�