XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150+^��,���/7�����T��8�箍l11i����[�Hkw�rpH��:�i�uG�������/)4�q��?#�����]�wX2���������׽�����e���{`���3_�[��UE��
AX��y�	�m�3�������f�E�ޯ97_���?�et@�7A>�G^���(3���Q��c�t�!�F `�sPя��Û}����}�u�[@���t�H�4�BX`ϋӿ߶�s���|
��8�	a�U�sxvC�=���
� ��0�r�C���h�w	�o�;�� q^ȡ�G'z��nZ����Q�,��)>���z�o��"_L��Rf*c�XlxV61EB     400      f0�ʄ`�:AS0bu���<�� ���I�A�������������_�z����� �/�5_������[���)M��dqZ�����az����IHLsw��F��J��i��4�dﹶ�({���g��g��W㶸0^�Ύ:��Z�-��hV(�rH��8b3�y7c�+��V+�᯽�HC��)�z�G{k��#���i?\�m㶎ü�sP��v�՛�����\6��n2����*�A�XlxV61EB     400     1a0@l�Lz��L�r��~�u�<�|1: t�[e[Pt��T���!y��3��h��Ǌ8���֦\�ȼf�#=���1z�c���9k8=2o���b�� �[~�b==G��q�l7l����F�#�~{��� �6W_^��/5��j���N���91X�gZ�u?��khGy~���TWP��f���	�%Q�˿��Od��5
'�0엍�Y�#��$a��P@�	<���'h���U����}s�(�gU�B&�k4��(q��zaz}�.�%6 ���C�V$�3��٤����)�z_ �lW���Qi���m�5�Y� ��+9}����v��#$˽���bi0��[o=���^R5B��.���ʸ�<">�.S��[��||'P<��]
�"��
G��yX��"Jo��$��XlxV61EB     400      f0G�Y�l�R](�'��1t�%P�/��ۉ��D�l骲�L�tI
�{ȨH��>��6�pe��BIV�"���\E�w�rP_z.K\�р~�i=���4����_����m'�	��E�z�N�&��6����J��|3; T��;��$@�q< W~􂋛nO���mWsM��#L!��+�o�g�衝Z��~4[g ��w�!��������R$^��l�b��mXlxV61EB     400     130���|V:���bݍ-/�<ԙ�j��+I=!�3�M+����|����k�R�U��4�Q�%����&w��;w�J�/pyA�d��_R��A� X$=EsV�r'�+��I�o�`I�,ƪC�M�ޖ>z�f-��P���ه�����@
d'1]��?�Q�A���6;����_3Ǜ��ڌ���Щ6��vȾ�Y� ��@g8_#��9<�)sǦlI��?�`%��D����
��8;��� �Q2��^� S8u����B��fdG����o*(d_+�@iyx� �A:rXlxV61EB     400     120����7����g��Jn}�  +]{�?}`���}�m9?j
Qﰮ��J�(��#r5FM��Ə��߀KI^g�ͫ���'x`��zvW�fphIu���:`�ė��XU����pV|}ƒ����]\rP��7�l�������෫/Ę
b��{�_�y�m�rm\`���cBIN�k��J\�C{s�N6���a��s�����Ո3�(mӳ���^��D?����NR��#4�S��nj�~.��js��V�2�Y�
����ue��(��U*�&���W��#)+�AXlxV61EB     400     100	9p��gQ'�{��U���
��,0U�U��J��NN�v]]�wbͷ.���W�Bu$���`͊|��O�T���x��JAI<�m`��ȧ��T9��,�%�],"�h�)�A!c��^�(��`���9��'d�\f�7c^�|퀬��6��JKl��@���*��z��ʡAWS\�� "(��ꄑ�|G���<�k1xY�{}��ҷ��q
S�f�tb"�OyWv{k�i���h��R���`�WXlxV61EB     400     160M��'�?k�`�����b��K>�������� FMuhk�o�t�\I2r�dhd���E�%b3���a��4��v��E�������|���':Ya�62K�V���ȉzxV���
�Z�����7�=G�'d�GLW��/��Z-�GDᏏ�g:f��V�
F?]��g��g\4e9f@�M�M&m�^7> ,?��*�bnݱ�bafU/Y3h�_�d�*^س���xz�E���P�j�GZUkҝ�%���ʙ��)�N
���Lu���U$Я��[W�B���
���t�]ɹz��$�jR������,O�f�
��L����.� W��V&��U��Um*�29Գ�5�2�h�]@XlxV61EB     400     160�_r��oC*�y  ��;e鼟@�"-��)��:	T�'4��G=�Q��X�ap�0�`k��<ʢ��'J���0�*БP��eY��;X9�֢��mr����u{~w��f��-'��A���X&���q1Xq��Ҷ�\2dѿ{�Q�E����&��7X��%����v��H:��8�PQ8.�w��Pu�� �fMb7�����~���>��)�_���Yk�t�m׽�i|��Yf\M�1p�Y}ͪ���/�-~	�����	X���PYѱ�Kت�������.�;��Ȓ�{��H�er��~�s��.�}:�~4��X]$$6�"	����]:��WXlxV61EB     400     1a0]{��R�1�+�n��2km�al� ZN2�D���g2J��c��'�#ď�l�)d�p�"%���1��/����C�UԌlֲ5!⋏�M�6��TŅi���WzhU�h��"�t�����ܮb���ܛ��t&���.t�k �ShY�(��j/��ܠ�����ȍy�
��A_�e�}W�0Twh��I���(~��{S�σ;�bt3���`\�O�<�4/#`��/��,�ouZyy�Q��(�^o{��*0M=ۧ:��H�b���K�O+��S��28t��o�l��wF�W�s�X�Fw�3�؍E��0��j2�I��m�j��ԍ]�Vz�g��<ZܦCmJi}D
� =���V��A�$% �z�#��  Z=�X�s^Y�&�4�m�U� �E��JPr=XhZ�L�Bޣ%�qXlxV61EB     400     160���}��^��6~5�CC���� 9�<�nKz�p��i�;�^^�8��n���fכ5���-�5w�yާ��6<�@g���&�h���󡣜�L������#��ﺯ)��|��Q�������Rˀ��h�d9/.v���G���Ť,��o3e�2獴ʈ��nE�9���Cd%b��U�&tGM�zA�w��|�e^�"�|�[��y.j��4J?�6���{�z�^��Z7�+e������M&G���`�� $K3��w1�!�;f�ד�Ի]%��e��2��ѹ�#!�@�qr���D͙i��)��6o�0n]�4(瑊+Ya�\�XlxV61EB     400     160�5od��b�V�	��t0p�\�J�d��J�%���:�8����z%l��m�3�R���]J���F{=��r�aW�\f�f��Ox���<r�f#Ό��ǒ���p\������=�PJ���m\��������)��� �$��hmR�P��,زw�^�b޸,���^��|	{�ՉY�K��M�]n�v�v}�|hr1iˬ?�D����Q��_#�)ew)��9�ձT��@��3y��8��ʡ�D·�1΃7��.��-ًL����G�a��Z �=�*e4���p���5[������@wF�E������
��O�z�>�H�g)2� K�[��+�8'��XlxV61EB     400     150��i#�G���e�S�3 PZ$��!�Ã�^�:i�d�n[�Q�d-3*�`����\m���_��A߯� d��ֶ'��i�ک�bN@jX/Q�%mش6c2�߹�?���,�9�0`#����y6�+[Xo��mʫ��"@ ���n�[P�Z�<c=귯�/8��y�ZR*����/�XsK��(kxZP�\1z,�8Ɣc�`;E�,J]���7�-cZ�褞�jިO7k�j�(�z(v�����m��)�8��n�z�ب�>�Vw��y�WV	�5� ��i��-RB�@ڡ`z�pt�昪5�w����=���7�����`�F�(	�t���u)\�.XlxV61EB     400     150��W�	,O�����4�3����M�A�����]L��l�m�ssF�����6yx]kp���+�<;�J�}�+�^\�r�'N^q_�|���Oj���=���b����H���}Dd�k��O�.mEX�?o(1��l( �ε��L��9v�<��7�r���cx��,�����PW�;of��I/�R:��L$ ��e(���`���vP�����})�!�U��eS�L���/�J��*P�&!�_\j�D~p)��H���h	��R���̕#��t�/	6�Rf��+�6eY�,��[�S�
��Rx��CZy���:�f�1�^5:�k|�Ӕ|�XlxV61EB     400     170�P	�3Ÿ;�d/�cݨ�7[)m����RQH�¬7�������H�D��5����Ks������ޜ!=���e��e�q՛�p0������)f9@.��Q q0g�L������w��ذ7�]�~9*��@蚦K�����c�ǦK
�*3)f���M �]��lgrd�P�Y/z���v����+ǅ��#zb�{fF�X��|6��ݣ7=h���&$�wKAN���q��$-w�yF�/�fԤ!�j|�)����Ͱ٪e��y��^!/~�4���Ix'�����v��L0!���%ԅSE���LK�'�c3��*o̿��g	J"ٓ������^8��c���I��Z��}�O�s��<�~�㨠�@�XlxV61EB     400     190��%^��6k���e��L�|�ۈ��-��|���p�V���52m�Wu-�����Ǯ�*��-C���k.��J3h!8���p�Y��];l�2i3�A�-}V���~
fv�sk{��X�eKS@Y��|�<��U�4������
���	�'k?�E�*�4��n[��JH�",��i���H��p�@�F�ˤv�@Ź�Lb l9�n|��k��$�ꍔ�t�L�Ҫ�I
L2�m?$����E�-^�T!����@y}[�ͱ��֨b���9h��	��Aڰ�`�	�Sᘳ�[-y���Mt��6��m[�X���wu�akp���?.��^�'4���:�Y*)��q�ת�d�.��ܺS4��=�.뢞��� �1F�e��0$��E���XlxV61EB     400     150w҅�Ǵ�6�[4PLg5���_����_�I��%Zy8�1����%�ՎO����6R��:�6�ª�Y�[G��cQ�P羨n%��S8��͌��f ]{$����E;���
�����g���%<0���fo��>�B���1�Dƒ屟��+�����t@9'�\�)�م㹨E����(TǵH�(�l�t�Z��?~��SO�-p�|ꐣ���"Ӄ>/��P3���S�ej*9Y��:�p���:�I�#�fϗ;���L�ڭ�T�5ֿ�u�Mr�[O�X����"c����z�Z�aX+�Z�8�$Z��r�|D����XlxV61EB     400     190��'��~w�r` u\�4F���>�&6�,���y�K#���c���<,����6��<������7�k�g�L�5��Yا�_k
ъ
��9̯��a�ɻGu,��P��y�$�}���^˃~�5�[m�f p����y��TH��u��B�1�kiIRp��Q%�7�����ڻr���yhe4�'q�T� � f�������rV0%	81���IÒ�P2.Q��eM�K�;�,��=&eÓ�������>��m�SF�/l��L(�R��ZW6�Vi	�9N0���ծ�V�b�$��u�����4X�|\CL��� �G�����d�퇊@u��~c�u�2V�u�|=������g��`'w�������I��TH�d3���0���9(��)���pXlxV61EB     400     1908Ӏ���e%�d7��80z��0x�!�&pHt��gNr�U[����a���x�u������ܘj�����l_�*���Z&TO|�v}����@{���Ic"Q{�\�ku���U*�'bq�w�xT��GU��Y�~ �f���+��e���3n��Z���Dh�I����!<O:T1~��+�Pl[��ƩY��v�ɿ�X��&o3����ƅG|>�H���4>�@�l��'�~��eg�$�,���l8�2�>#�f����K�#��չ U>�� ��uYq�w���{7�C*��l����W[�qh2g�3���lÃ���� F�ؚ���5��<N���b΃�Z&w��;�*�j���Ϥ�}K�^Q2.�+�qTz�>��M�5c":XlxV61EB     400     170��~9NV:�+F�����)��T���#/��W�F�: ��bI�f�^��6��X�|c�/�Ls��������n!���S���<�%.����CY��G���>���u�_��U~�ƽz�Kt��͍��(-t�B}�\6`'C����9z��Ҏ�YBG.��@e�g�ԇ��v[5�+��N���hq�Z*t_	|���u��"7��Q�$+_M�dS�+.~d1.���L����n�ςR=LnL���\1����49L�'y�N��D���7���C&�tũ�T�ʞ�2B-<׫~�j7^w�_����AF"c|�Z�� �7F[��F�8//�-#�z3��s�a�{���x8ĦS/�ddćZXlxV61EB     400     180.#� ؤ���i���z3SI ��TGg�?���8q�8�$���E�AՖ�4�.�1)� 5`:��\Vx>�Y�30��M�s2�?�UwJ����c�b��ͅ�OHtEEz��X缪����(�Q�������$6ʂ��!�f.��z۫���}�
�Uo�]4�;�壇�wy����)�c��T�Q���'?]ҫ�:�K�Zk�O�Hh�����RdM5��=<k@�<���E/�R��Q�{�*�A���6-0������p��'?��Ĩ�J@Y?��ʚO6��,*�P�0	�s�x���e��M�����w�����C�I�BW��19���q���T%7?_���j��kZ*�.�"����2֑��XlxV61EB     400     180���� �~�}~��I-�9��g�w"n�I���3[z�Ρ�݋'Օz�,�֘�0n@��*\��O�,=X�&@{�i�ad/���G\�P
}��Gs����.z���ERԩ� �z�����ȹJ}��a�~��?ھ̚�����N�{AM�ӻ�H����]Y�|������ .��K�V�i�H!*�+b:�S��k=&�z	;Չ�C�ܪ�k��,���+
{X$0��cn� �V���'�V�bO��"`�H�B� \���B0�G�H��氉R�̜il��"����7.�E���6ؽ{c��p9�>����7$,V5J�M1��u�wN�E��r��^�a�����|)� y��Q�Y�T�[�Q�{�$�����d7XlxV61EB     400     120%r~�&����ʩ�p����\Z�YM_Ĝ���q4_���B��I
\�F^�~])Kd�a�Z9�r9d�+��z��V��|Sb�aςQ���h;S��6��"�?� ���,`"v����=��mh������!�\���H��?��U�����I�ƞFd�����Gͯ::�j�����9^N���u�ɣor �>GQw�&i��&:�L�R��r��V��7\�s?I�!AO�pk���}�0"�L�M�1�<%��� j�Tgѯ�kT�?a�w�\��+�f���ׁA~XlxV61EB     400     160,+uMw��"?X��D����QՆnv�ZQ⮈흷��S3L�' �O%�bѨ�d[�m�)}BZP�F5�e�;�EY_�=�*��mR'����6��#m��L�٧!�s��c�S�J�ϓZ��>��^�����IwvZ�l}b�9����s�B�ݳy��΄=��[�j��o�g���o��J�=���¦���O"�7�L���n�j���Y!��Iڧ�����={'�$`�kF�j�j������t I0�j1��g��%�t:��E��R���:��8|�*���~G`��#�H�g����j�����.��["��(�0Y�J���v�h	�|�W�؊XlxV61EB     400     120�+uǎG���X4rb�"H��ٰ �S-�>t~�yN>Hj>3%�_�4�g�F~����X��1�Ĉ�D�L�|�\��O�-�Q�P�F������n��&��՜ddA��d�V;|ƿHN/hj�J��-�_3�)���<��U-��޹3��8ˊu�	T�Q4.�< �*��Q'�͟]��Nf�j��{8��!,��O&��d�<�Uok�p���`'�{~Ж&.J��^Z�1f�>h#���'�K��� KH��-�: ���	PE"�xK%�8MDY�FXlxV61EB     400     160:��L��٦�j�N�<��(�JU���<'3����5}�G!��!�o�h#>ǩː����yQo{��.�U�M��B�)GiZP��צ�"�;\-��b�+�bb��+m.����%��A��Y�^%W�0$Ba�vGF搎�e��·D�~��SDe����u���+��b���݊Q��~��y���!0�mo!62��y�ش�q�y��?aĆ��MW�d�L�+���-�I���c�zZR����g�5�y\=Ev6��bA�\P�5(���?���F�☏l�`m]�qz���jX���/�
����5ێ�M����	-H���U���+�Mge�	cXlxV61EB     400     190� �U^����s�,���CP�Hs��Q��9���.�1�́r;*�^�NZ�I=S�&��7ܿ��Ի�q��F�ɻտJ�s�U��#���V����@���X=p���erH������fG.'��Wnӥ�\��5D޴�(}{���W�OC�"�#��'֯�=�=�"��\�(SK�kй��ݽ��IY����7AZĲ5����3��v,��ឯ��J1� ��M��Ä��e���Gw ;�`�t*�����{X�z;''�=�S��h�UYC�wzk[�j�ܹC喛I����>�j����nB�}G�6���Ƹ^Lŗvs��gi)Z�lB���m�f^�����E�l-��o+����i�j��]�#}�WT4[*X!�4H�{���*�_v$�F�V�XlxV61EB     400     120�hh�Z�?I74�	�Mr�_�	��0��=�L��u��>�p��hR��Zp�o<)��8:yQ8��E� ��;(�ѩJ�m�����YP��X��o�X��<S���c��׈��J^��Wƍ}���TY�í����+@ {@Y�=������S�]�(f{D�tI���W]�4�	wn����=@�3Oi�t�A	WQ�@����I�{D�}���ܝO�&���%RrPFˑ)O'/����W��Yr$�Rݶ�hi�Ysy�3���m18r��_'�3y����f��XlxV61EB     400     160�]�[��I+Z�x�� �	m�eZ��Jz�;�'G���a�k�!*`Ώf��������������G^��EK�6E�愪�4T�/eS�F�����e�#`<W��!~�$e�MW}��l�� ���56�R���Uƃ�m�d+э�G��{1,� �Ǌ,�m�eLފ�1�|	g6��4y����A�՗춭��՛�����ab?�b���P�	�1Z��r@�2p�y�82�&R��6Gg�bn��M�;ދi��ׯ�ia6��M�����-]�ɿ����q�sTBD|�$��th����zR�m���j�4�n�h Խ�Zy��>`���t}h?9;lQeX�I��k�XlxV61EB     400     120��Y=��%v�9U �l��n����d�{��]]�9�u:��G�4ʖA:'J�Bz�%�yf`$��Ua���>~���[���#:�*N}s����4x�yMR�w�OC���}����%�����r4]����g�s�O�0!�`v���ʭ�{]�1�e�/ˎG{$�I��;�F�,�=�@.H���;���5���4��U2Y�m7�29+7�R�����!1.o�d�o�y�Z����
D�K&�R�9(5�t���)��қ& �z��4��q��1yXlxV61EB     400     130`;��)���B�8�7���+΅�e�ν0-)�r������K�v�B͐��Qj�[e��&c�VBR%!�ܩ�5�i.�.�*�9���ڶ�#_�O�8�潷E�cWOyyLt�
�b���`"�(u��B1V�k��,yt�zB��J�����H�������f��1ՊIw�q΃V�H�Kn��.�G�^���
�ln�4�3������|��'K�|ׁ��h��4jn���UV��,�ԡ�L1�%�uT�
�Mg|_&0,b��̊��E5�&ޘs����ɰ�E^�ۘ���KXlxV61EB     307     100�p����b%��~sEyѺ�mIN����>�U�d��a||x�~G42�L���p�icG��3���L���1k��������^�N�r�E���vf�m�������������j�F�AQi��9)�Bÿ� 0���~h�CC���S�(�Y�@��*O��*4��е�H���u�E� �e�z+=U2"� I�)~�`� v�u���Q�=�X��3O.�������,�!�م����Ej���