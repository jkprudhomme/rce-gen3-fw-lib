XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180+4[�@�+]��3d[�4�c���R�;��/�M0 ��뭜di`���/2�;5�J����N
��f9�\k�����x��fuҪ��PYW�ճ9?r#�cIg�=�Z���bC'-�5*x�x�[�)����a���;UHh��K�u�Y��ˬ����$��I���$��i��8(�M��P0׎��d4�����oo^�:r�L��[P�](v��8�����Ц�M�le4��?�n��K���9бZ�+�3Sw����*��W���]��>��L�q"q���Y���T��k�h�>L�.�s@���.�N����޺��0��]'r#��ᕖ���t��=��U34yɀ�ԯ�,CO��|g�}��c0�g�6�~�u<+�Ԓi�XlxV61EB     400     120u����WH��h�Fz��gƞc D�rE�����)���iw�m6���$4��λ/�7�U@�p��ޥ#)*�u <o��7�)��[1�����g�Z�:�Yr3�8fE�x�@��p�$�K��i�̷=p%���a�ɨ�q��m\����x���M�qQ�<�$��kCx�/03v0�iG�ߨ��Y��Թ4j+
�o a;_ׂ�n��]�lPqiڍ��2����CG�f�Njؒ�#e+��A�1�0�m�"$=��P/�������fKè���3�b�T�#��dj\H�XlxV61EB     400     110��E���~v�Y���_�ңO�B[A=j�L{@KQ.oHXYޱ$`\��@�������>c�]@#�8��gt�U�/���B���:'%�Y�'x��f�.��/P��NSǸ#�My��)�����E�P&���W�I��g}P!�7p-P��8�&��7W�P�¼QB2�k���@�G���n)	k�M(o���"
/�VM�.���錊#�6����)���.*E�.J���*��ڊ��l�S��Nt�3K�7����
O��Xk���O�TXlxV61EB     400     110�5cK�������M���E��w#�-�,-M��9\�0rK�V_5YN�#��o�/��M�H|��;�\yY��I�g��Bה4����;��3��z�<k ��3B��I���W��[��\9J!ފ��T:���D��Ŭ�{�$Am	/z��h����8t�w����
�Ȏp2�� �۰d����p���6��=e��&�Ia|�ƞo��3�Lܐ,+�vWW�7�
�5)�w�q3Z�K��ip�͇h�MCΈ>d�tXlxV61EB     400      e0\�͒`��as�C�'����_���/��)��N��(%��bb�uD�C-�u�kO�yZZ�5�lQx�!��
���Z�
'�t��i�]d׆�F�8_�$U�K=�jɟ�RŢBf�c|(�c0A����B���)��Ji,ih�M\Q��qF#W#��3�V�׭��l�"�ۙ`���'�&=Li6wF�ڴ]�FV2��ׇ��\�ܛ����9ĴXlxV61EB     400      e0�"��.�%�9�Љ{�
A
qUW^N�J�b�s��nH(�׸ªp� ~�a-��}yr��ޟ��uy�Am{�<F�E���禰�0�P��N�)�����Os)Qb�X|_�+�5�py�{��3�� 0��zj}�}�g�Zq� �|'-���r)�,Ζ9ruS�Ħ��8�I5��Hݏ&Ȃ�+"�3�!ݐֹ!-o��9�kb�a"�}���/S+�XlxV61EB     400      f0p��FKS����U���͠�O�%�>�&ހ��ت!�N����[.�A����)�x�Ϣ�_ 2o)��O��.�}.��M�;j�5܏.���_�,9cj��Di@[6�`�$��IK���8���q��]?).�8��P�~�Vw�<4�LE��z��c�n-K�[3W䓪E�͑��L�oE<yD�<T����*�-���-�ζ !�W�H r�Z����G��+ͤ�6p}bI�=ɡ.{�+�XlxV61EB     400     1a0Ǩ��k���%ޑ�8 �Rw���=7�'�6-�6��¦�C�&s�u/�V��L9�194Ǣ�x�I�d�w92������t�^�,�qu���Ek�ٓL�j-�SQ{�N�ޡ��U`򼆰�X�j�;Bh��9O��%`y�@��c3�.GUU���\�����m�۝aL�}�v��!�Az��:`�=1��=���v�m���)�Zn"��y���\��@Y� �+�nǎ�
\"�J�P��Se�v���k���O��A_�����f	Ej���壥��+�� ���s#f;�����C�F�>��6 �7i�	���H�u3���wOI���ck���#܉{�E��� E�6��S�(��*�����y*�^���$�Bђ�o̟����Y��(1<=�e"y�'���XlxV61EB     400     150�*����+�Κ���Hh9Dg�)J�==��N�+G�g��ǞF��4RA�Uzlv�ݹ����I���D�l��k�.�Ȉ�{�i{/?+�,W[�
6��}����/ m�,�Jص&�Г�3��Qs4���8�YW�`�\�Λ�G-��ݝB̨ ��N��h�׈2�t�����W�s3�Uʭ��P��KX�i2���8�[��'��y�cO�׾��N$�����-�\o���x���&���h�k��*ɢ�]tL�r�Ï�%��
Ч;�3�HϷ말��(�E�P!�e��r����J���U:`��tu?��5o�MԻ|ۋ�R�=tu$XlxV61EB     400     110�u�*�Oz��{Z-ޙ���gy��񤈍#���:%�Wb|�K�\�~?�~�ZűN:/���UU[vpmԐ=�L��$�6���m��ZX�����ޏIH4H2(WGx�$��	�ތn�i�]��A�}("��.%�s����_W���0�#�(�҆L~y�H�pP&�9�������+lk;:-�����]7��,'0�(���%��@$B Q�g/e%݀T�6�e~,�"����KoP�QTz(�p���M&K��#4JF���N�XlxV61EB     400     150�i�x���٥Κ��?�vY��Ż}a}�BPsт��!�Vܘ!Qދ�z�t�(]�:��+Xg�����k�u9SI��蹁��5�_�.��T���e�^S�gg4֞a0�����F���s>��:�G�,�@��+��[���@�#K���]�<m�'�����S���Pd�+�x�i}f�k4�<z:@��C��.V3{@v,�+@Fw�A"|���®��)�L�&?�{�>�I�$LN%P��o\-�]��4@�L�Ȼ�8�^��^xE/uh�L���&hC@�-1�~"�1��R'�=�eF&T�iu	��Ƞ;��較����|׺v��ʬ�w*XlxV61EB     400     110x�������>���K]fςde<���q��6�ska�!�J�8�����*�s�b�B?��R�t�'̯�HG����M�KX	��w���)dI�{AҀ?��װ��b�9�������$��I3v���8�3[`��8���>ML�O-�-k�T��,������Z���s��9��'w�E%�Ѱo�y[h�ю��� �&����o?7��oi�V��h�J��� [��3���a�-��b��eñb4`T�@�X 4�Β���XlxV61EB     400     140��)A_���ɑGsֽ��[�[bkU�"�b�.���'��a�z��}q{���~n߰l*3�+;<#0���) Un��^�5J�Ȁ���R��+y�b�L�HPl��<^�V�� ���Hk.��T.G�0�`m/�ϲGp��ِ����Ul�t��;����%}d�T؉PD�yܣU���F��>!��{V]�-OI-�#f}�5Q)��)ꨎ�,k�7�A� �l<��@����^f�y�$�u��f髜iըfBQ�l�5�L2���e!�:�Xt�ɛ��㌋[���6�V�o�tP�6^V�$����y֑z� /�XlxV61EB     400     110�yQ$��iiˇ�%��?��Z����:V3J"�g�~�)=�ʡ����qHuXq'�t�6������]���=gI���$�w���{��lI�U�8\ҬC☇Q,��ߜZ�V�aۧ��b=�2��)'���%}�5X�G�>|���rJ���'��
�Ӏ��Ͷ�))� ֠��'\�f��'�r��'����`�R��r���������:]���Lv=��: ���e>]Y;E���7��_Ot	����6���)�¤��"����XlxV61EB     400      e0C���5��p�)
ޠ/����0��G:6v��� ԙ��]��_:p6�,y�|O�G,GG��B��u,] .�a~��N(��+�,����D_y����X�eծ��X�RR�p�c(7M��oA��1���fDJN�s5���m���#E|��pj)s�zG`]�ɨ�o�~޺$;%�ު�9HΩ�,Rf&��'a@�(���g�N�Y�Q��^�^�oh�XlxV61EB     400     170����]�� � ��&������3Z��?�8*�#s����cC5�hq��^0�;�����yَ���<�[��7�m�����@��w	�"�lҫ�:Ђ��kT\��#�x���2����;SG�qs��S�n�Oh9V�e<T�S���_a�1޽A�#i=�k�v�cR�뎱���O��E^�)���s��DO�po��w�lc�ryI������Yhߍ�*6�eM��ـa�&
��h�Ds�,
�Ex���m�qΊ�-ʭ]��|��V�8�d�ۙݚgDQ��l�y�~�� �)e�MnQw����׿�騠��KH��4@츰�ç!���!�9>XrPw=t�r�;O:��Qm1C��3��XlxV61EB     400      d0'
�[~���i��t�-�e��]��UT������ҳ�t܅��b�S5H�A�&�_�n���zV�2_�˔?���s伓D���\��+1S�@�-.�=� \�w��H �N�/$K��Z�������?�rK/fi�c N�f���"%5�#��\�h�o�v�S��gF�#�8S�o���֥�}Sx����/3��nVI� �^�� Y�iXlxV61EB     400     110S��sZ#-ߪ�_�\�vd��Q#r���{/�X~W+��հj�|�ϫR�>tI��������  �d7mB�|���,dk9#%]���1� ��� {a��C�b�voє�1o4��r/[��t+�B5��Z"�Y�ت���<�j:��՞d���0�g�%0��s��;��I��w��k��­#b�[H�[]6.L�E�C-Nˈ���2/ᮨ+�)S&�h�����e��\��)��Ŧ�|�#q�ޟ9?�l��ip�IXlxV61EB     400      b0�r�\��������?QRQ�r����q�EfF��Aϔh3���֩���s�ݤ�e�dP��+̇��z9n.0���Aj�tP��o uJ�w ��D����J�\��'�ى�*�(No�ã��[+��]{��>f��dH�2�F�7ծP�����J[m�n�ү�>���*�a��"��,�XlxV61EB     400     100|�/��M�+G!��H��j�"�{�8�>E�v���S���ŝ �!�w�//��dT�,��J�E��%Û���u����֑�'�m�!YA�޶���[�LdX�K�>��`��)+Tk���Pq��Rdܒ�k����S��ҤU~�~�2դ���
���`*����(��k�+�kج�H*�7�
㌣#�!R��HJ���$�C@�B�엇�7�U��� ��>�ő�j�J7���Ƙ�q\6H4�{�� zS��XlxV61EB     400      d0�\4y<j$�q7����c�Q]Sb��z��?ؿ�҉�+-0�z�-��\�A�zc{�4��g'ۥ��[0VoU�eiaK�6��c����������U����s�[�����t�b�Hnȭpz-U*�.��c����c��&�X��;��$��=���IBɗI8�vv|{NɞK�����}���u�~:;!����¡�&4 x5�,�XlxV61EB     400     110Ă��t-~�xFRɹ�
��{�J5��Դ��s�lM�+��C��r�8�L�1�C�y�`Ћ�.�u�����o	�wj*3��A�d�dYQ���ʮ�O��wU\�< P�-EF�]_�G֯�[t�>==cj�W7�C��ТI�BQ���3rflO\��� mq������2�@5-G��]�v�6���Z
E��K'X������<��25�Ae���=�{�� ��"�&�:���]���n��R:-I����7��͗�}G,��-؈�֟�XlxV61EB     400     190p��l�GZ��ϡ�I�2g26���T��e����g+�6l��E�����Ξe��M�A��^�f]�L������������"-,C�Βq�
���4a��G�7��x�!ȏ�nB</q�]��+�/��["����S��Z��gV���):�6#�W�/z��&|�=9e�̭�S-rB�r���r���?�@r����DEy�F����է�V~$�sK�� 4r�T�{��F��gcv�A�i�?E��>n�l&30�6�`	2H��{�Ɗ|�;�?�^?����D����j��&bu�Y��(��f2q:�"��>qn' ��	�L<,����z����$HJ�}VR�C��p՟u��pdb7M����ڷ:��w���ZY��Y�����6���\��<�V���6XlxV61EB     400     1a0;���S�M6��g�t�u�X
�.gg�$��&��}6p:'z��c���^D�{_A@(i{�[�*x��m��˖ϫ̔a̛�kK��i�2̃�B��Ik��k�V�\��
��=H�L�h��uS�����py���uď����K�23��C��\�=��.��~^x�E����������.BsmN�e��Y,�i�|�$�3u��VN��é�A⡬�Lg�Ë_<7������i_��֌�@00���C�F[�q����>�]>zBY�[���m��O
���2��P�ҔTo��yipMg,���!蝃wlJ&�0��j�d�Y6�q��6�YPڶ�%wH7/��W���1"���6�	ʢͿ�~��#�VO��P�<&�/��0Yb>��ʺ^YfS�)~�!cpXlxV61EB     400     190(��^C�P��^� 
��� ˜�7��.@ͯem��@Q��
��4�Co��["������|��!��h3�}H��[D'�ab�Rm�M��Oe�����6�c���w�����G���?�h󗍙H���~[Z?͋*�w���?�ĤK\�+q�WC)��4\����o��>�5��Q��B����Ȗ��K@��)�:;0	��̹���Cd-�]A.re�f�9Y�f�tL苎B�DN���2H=�6zMv���2S��ڸ���&�v�Yr`���N�U�(8�΀�y�-('��5���,.�JI@&X�D{#U�,{뾅H�M(m��	��f��r����Q�{����m�l�˫�v~*<C�[�U�X��]�ѐ�����eg��LnyABXlxV61EB     400     180M�;ܒ/$YP�}t�}L��� Ts��e��R�PW��֬pu�8қX�D7;����=��L���B��0���/��x�@6|cX7:-M�(Hy��/U��r(S,t�DL3y�=��q@ٛ4�hHtB8-��|����D�x4���i���О������q?:~$)~����(d�*\ʎQ,	V��{�9�ډa�q�[&�~a|B_�� ������tF"̈N!���L������!͜�^W^o�}k��5�bҹ }��%��3S���bJ������x��g�n�*��p����x�n������JP�u6a(���@��q�@S�G~'̾`�j5�o��U$J�.�tCP�7�k��.�=�2XlxV61EB     400     190QL��Њ�d�m;��X-7�*H��6}/���b��-��Q��^N1��"afy�ܸ�^(5�vŌY��*����]��/��������Bw��bf�xWn��ŏc�ft���]`�ē&�������hQk�w���c�7�=�w���˭zT��m�戜Y�=��������|XlG��>k��
J��`	��80ڍ)�XNM�=Q��t݋���k���W+-) ԰�4�&V��aä��B�3IS���s�X��UhO��;�7�⦘H�l���S�O��)��6�d
�V��e�&�z��z3�D����nta��f��Rs���U��hsD���#�ܒBK����xդ.�B&e^��%+��>Ǿ1j�{/���oJB���O�+��F��K���~�Cj�XlxV61EB     400     1a0�ʩS���H�uoY��?�}�I@Ǭ�:�c��3q�kUt�ٝ>�,FRo� t���:-rv�����Hx>S߹��%��G��������P�i5���mSN��h��q�'	�d��
"	�Ij苦�K!ټ��D��ڰ��t=�/�c�ڳ��g�6��lxU��h�ù���H$�����ƁK_q�TM�v;���� A���17Ϟ���#�}�p��[�ubh�r{:���n�0|�`І�/��[�:R*؄����(vn`��^�7tW���B�h��q�D����Ñ/��Ķ���T��D�!^C������9-��H�['��W�g�8�-ܪ՜h�S��v�b��aP�5�!�~Єh2�YG`pJT@��e��5��""T�,3HNO�GV��r�j��K���*����</��	�_qXlxV61EB     400     190ġ������+
Q��t�n�aӗ�#S�
�ro-b��\{U�P!�?�->��P�u]0�7����P��Tf\&����o��u�;R`��۟:���S�we�o��Y>�WJvٝQ�|؈4��Vz�b�,mg�Okԁ�Q����j��Pg2���>��������u+�=����*��{\r$�S��L�A��A:��=ʖ�NA����T	] ���p��~K�Ph��.�)���Ot�!�FDܩC, j!�B��7�S�v6;gW��w���	��4z�G�2<I���؉�n��� 7���ɚ�-Izr����m�x���T�o(��T�yY�n�g�1�7���hCl�`ے��9^��ýV���%Yc
U@���wO���4��Y)tA �[��؝�XlxV61EB     400     100�#��υ~u�H�R:R�����B�۝�e����d��q)H8�$	������U��v��i�ı���"�d;����4����� ��p0u�=���(�Ӿ���8v;;:� �P�����@.���3O��N���� Qy�=�(v��0J{c�ύ�'Wj�H__ML�Mfz�$�� m�,���6JԜ��9�ә��.�,���8NA��u6��nnI^ݭKx�� ��lu�*��VS�q����wXlxV61EB     400     1a0ʈc�S�}"�rX��RfG�u�/�H>��I������yM�Q4w�ԉ30Xo���`͸�$�i��W�KI�:9�dV6<!�b��d��Cg/ԭ�AK=��	ŬxF�-J\�ũT�Շ4���.�<����q�v0�0�A����SdN�QȞ�:b��2M���\��ٻ/�Y�n�..xX}�Ov���/vv��-YF� C����M�B��(���w��h��㡒�*y�O�lɁs��u���3��� ���$��-��)��S���~�l�����<� 9#اm���ބe�f:`�"�=V�]��F�ڳ�L4�kX��Ѷ�vU�����V�\��+�Y�Q��L���a�*sٳ��q(��.ON�>�A�o�n��FR�����A��z����5}U]���XlxV61EB     400     170��Ȉh9��S�Ș�K:}�c'1��r��+�[��G�A�ћ���q��v�t/Lwh�r�2ߖ,��y�g�i���L�`���2�
� /���.�{�뷎y~n��JBO�*�XǑ��J-SK�� -�*^���z�r���(-M
���㓪)�)�Tg;h��#h֡��i-�鷜r�I�0p��}Ź�G6�2@�v�b2NK�n;�"H�D�_�[���5���N���]��b�_�ӦQT���3?$��{+����頞/�z>��)@����n�?M�r�6Eg_��
4�K���ެ��+���\����Nnơ�,��fe�(.�f�aí)���!r�L�9�FEG�_|DD��db�X���XlxV61EB     400     1a0O�%��0��?�� AL��erõ���-M�e�ǰaˣ��+	���<���2M� �����6��������K��}�.k��Yn`&���t4:b�־S��7Ý���e��ۧ{�Ǧ�\�LR�ޕ�D��G�q0�x-%��s�����^����#w�PS��]!�|i?�B� �S8�'��vL�>'X(�/�����f�2�_�gxl�Ϩ!+�ptI�c_�q,��S��T��2��������ig:B�����V?�jaᇾ� ]���G�`[~��T�'���W�s��i3=d�Ҏ�m��oj�ٓk:�Ӵ����z��k�Z=�4:�O5��	���tux����\��ƒ ���� O��3�\�m�Oմ�_�ztf�#�%���v�V)��XlxV61EB     400     1a0t6wI�~sf�\�z1k �x)����LkEhQ�W�It����44*t�����d��~���ޫ�.�c��2/�����m����D&�x�П����\gd*.�$�Ud���,*⅖����3HqJ�Y����!'���hbY�"��2tLݦfl�YM\�v#ҿ�!�/7��T�-u8�n��L�2'�<zH���=�U:�k�u �?�����W��?���@���G#G�$^�D<�d�i�(���%�ghc��r�O<:Gu����Ʋq�]F��Gɿ����ߨ�$?*@��X�8i����!���}p.���J<�������4y�I״���L]]�=��&��<)�k�PsB>&�k@���A���j����(�{�Zs��V4\5Z�c�
��}�t��)<�XlxV61EB     400     150��OG�)rxt&�G@���7�3s�� AO�ۦ2FKiu��Eۼ;5�Mq��,�[���O��
�G�#�'�~��&�~z]H���Kco`f��tL�c��`��P����أ9�{��D���6�N:
����j���*;X�M�ы��)�N��nz;�O|(}0p�B$	�o�i���6�{9s���'�vu�+�^��`��D�v5�u�`�r�!C��(�;�
��2E�>nT1�k����2J1�	���!xk8������䞝��3I����Rٻ3kV�T��2�u@n!I@�Cv����-cч���)x�i��)y�A^�XlxV61EB     400     190D��-I���tS��Mm��|~u��~6�܁P�bp�xigW/�>����e�n�p:��t�\.<���NʻI�S1�Rf���=!tݾD?y�&+�#��@�	kΟlDܹ�+	����jI�zL���̗�^ҍ.P��'wcOx���x��4��� ���}/G8!K5Ʒϋg�����u)��r�,�3��>[b��7�j�vAR�2z[��Z6�_���N����,�9�D��C{��ra�r%�U���eg1HxqI���ߘJj]�Q\�~	+���Qɺ�)��B�2I��=�Wi�m `�)� 
��%�<��������cnl��SY��H�">�a�����,�_����w7P@�����5qnҧP��pv�S�۴۾��H�{��0�_���gXlxV61EB     400     190�씉�V�&#I�l�����[�������gP��B*+��)��ݰ�pV��D�vw��WD1�"Hm��a�g���yqk0�Ѩx�z%��?1f85/�k�mJAr�������q��kĿ�[o돨"!���cka4@�@��5�}>4�l0?l�4�'4*������Y~��t��� �;�3�y{ye���>��	"�r�~u�QqGY~�zZ�1Ƴ]2����=�\<�jmV <5�!V:��9@4�p{���|�;��8	�	ar�&l#u�!f�Y��� 5�ԬAB.3�VN�̪�_����w�[�/0�+��/���\��r���AV��~c�h�_�O�8$��|�]�y&U#���D���^���;?��K�覆��0��&�r1�XlxV61EB     400     190-f�*=
�🺷�� ΞE�b+�+hO��y�+��#%W8?�8VM�[�-�k�����}������mY̚��:>Q�tm�Z��[�"�c��� �=�J|�Ez�xd	U�V�uNl�j;���d~��<�n�_
߮�Q�I
4Q������1;گ�����a��S\��O�+z�"�p��nú�&a�Y������#�-*�_�)�"�N9iv��%������5fgQ >;	��h��b��1Ɍ{<����_�R���d�P� ��=kwB�)M��E�������w�;��oֲآ�V���{l��w��B��,S�n�6󑊙�O�k�(�,�CA&I?�)�w��������,��^��NI�m�o���L��8�$��r0��4�XlxV61EB     400     100]��Ȭ/-]��7QNe�+���}ر�b�m�����tZ���WZ�B�<_�Q�_�E�X�Փ�	7�'�������O����\~��8�<>�j��'`�i�??X�_)+Gnw�Ck�c����	\8kv��������R�<U5Rax7+�Y3F!���/�#�w�h��?s̀ X���X��3W??C��U�Ǥ�(!��ŧ����qs����`C%ge������/F�V%��Ǥ������[w"�qoXlxV61EB     400     160�a<*r� �+� �|l%t�r����$�zcL��� ����7^� ���z�]@y�?>tA�1T-�!�}!7�|�f;%�7�>��i���|�\2���hE8b���`R���l���b���H�ѕ�����:�%l���A����9��$�!�C��R�E^%u����E3	�n/�ҝ����ƺ#��#��k���A�qX�­�� l�5�!�w��OS�����U9��i���ď���9������� ��y�������«���=�q������V"qb-گD]$��l�����1m�����$�������;}���c0:ܙ�֜P���XlxV61EB     400     140}\5��Z�_�<h,��Y���ɛ|�A/v T�0�#3���J�iJ	&)����y�\�����OSٿ|@%O#P�9c�c��1�<sv�jczr�1�w����צ'�)߇q�51�0�T^���:���~�@?@��cD��y��̔��Q|��Aϰ�[,�r�f�E��o|���iw�I��Y��#:	a�|�[q��t� D��г���Nݜ���8�7��s��tEߒ�����Բ@���,iR�����m=����Y̛]��i�R?a�<F��w{7�9Y����%"9�]��B�8�5V��t�"b	XlxV61EB     400     150��EP�6�tf�.��>Kd�3�`ZJ�:�B϶��Q�R��������͈�����H~�R�0�s9gV���K��R���J�d~�%}��CI�]7-�A/��_5n[�e�31�W_h��I~��밄��
��J1�ӌC�6	%7��_9��('O�X3B��Z[�F�e�RH�G����p��?�3;�$���JD�ڟDK�Z�^�Fa~涆�GǙ�e����~���ԁ%G���x�s��J��Ra�I�>����x7nl�%0�d��ܣ�T��<Y]�xR2xXϞ��̊��z��8�$��D�b�h���`$[��[[2������N���5��iiXlxV61EB     400     160��=mn���ڙ�ğڠ��P5 I��3�O{����R��lRY���YT���������D�3������6�݀]ټ�Yl��	��/����^��)"ϵ٫��P�if0�ΈJ�E-,.������W��X"R�s�I�@^�끨<���?�'�%�,�Y�l-X���Y��$�*	�����rs4P�G�ñ�+˥�F�Fm��g�L��[��PSW�hO�ˮ�"As�y�d��%�NN/�`4����<$�� ��TS]}�SF�����|�8nD ��,�O[�5�;KOOȔq�� p�v�%�ߎ��{k�E����/��p�Ö��]�e���M6�r��XlxV61EB     400     140�����Ѫ��ڀ/-;��a�j�5�����P���;�u>�X�x�q�^���u�F�1��dt��#��L_y�"�,�e0�CCYgJf��:7�QE��PZ{�P�- �� �8��ja�e����k�����[�/�Bn�M����U'�=k(0Ɗm�}���2�ǫ֨EȞG�_����G�CZ-�s���Е�+��-�ٓ��`�n��L����4AG{�c��]���x�SF.G[����+�駡���5�SD=��ԟUyT�>k�`�Ltω:e��H�p/�T'�?5�4!�{��[�OW�%Lf�	���ڐ�&XlxV61EB     400     130��ԁ��j�麌U��bJ	�A�%�VB��kc2sB0�?�ZF۩;���M"�h�g� �0�0�͌�!��Y��z�7�ɡ�Q$EV%���06�85�d`f�g���W���Bџ�b+;�8��z$c�<E��D]�1�S*B��Zz�5���Gy�)D(�⑕.�.W��)9�B��XzM0���9u�*r!}�q/e=z��`�V��2�)��-�c$dL�OL�l�֨G΋�z�Z;,q�=��@�B�)��#�����T�؉.vw|*�Wݐ�Oa�r�������d�Q��77�n3,vXlxV61EB     400     1b0"�̓��M�>�k�}f�Gh#P+(C�*ɏ�ߚ�C�yF��-�vϰ�9� o�V�N)C7��:F�=j�0X��I�3T�Ȱ��5& �7� ϔ�HMx�$|(/�|p}JL+�W�z�U��^e�R4ԞްBR-��� �� ���X��f=w>=�0bR/�&�p�Z���)8�;@�ǩ�	�Z�b£|���\Пl ��@���G����!�!᲼6�-�
���f)D*�~��;6���}M�^����,�e?EqSe �u0�*�������NY�M/��S����fxħ�%���R�x���.~&�<
��9j|6Bfe����E�����#��2S����<x(�O�HI������W��m.���Xm2���"��\=H��ې�&b$����lj�C��GϽ.�s���y�s0m�o�`XlxV61EB     400     160�I��˲1 .���IӶ����dOq$y˚<�����Ac��-_�;����+!�	�]��`��	,���S�g�5����e�5�f�q�E�&��l� �� SR�?&FH�Oa�?�e`�,�5��?��B���j}G�gB��C-Y���>a���<J�ޚ�餛�+�I�:�� �*�����'�o,J7��_d��K� ņ� "G�u�M<l��5] 	U��^&�a�31��!W~�����2=��T��(����m�7oN$����;�~&��R"��xC�uG3sT�!�a���X^��o��qhA��X��x�2�u��w��|����{ɲ<�����`ЧXlxV61EB     400     190��5QH���B�~ˡ0NC۰��Z& K��?	ੈII.�(�2�y��婻|�5��Q�rJ�AhX�"1��C�r1}����+��D��E�M�`�Ҳ��B@��'��AfA�ϻR"
�@������p(��vǌ������dh#}��/��iH]�E�a��_ �oܣ�7��7���Ŧ�x sdc�6.yȣ�kG�l9�B�/Q��Ĥg�~E�����`��]���Ш��"������Q��r���ֶ� �p�{����.�ӄ�w>ę(e�æQa��FQmi�-��'�,Kf�P���>�e����GW�_�v���X��=��0���J��8�q�3F`�:Ђg�KM7�^I��mˍ���jJq�8�r��:�z�)��P �=�r�XlxV61EB     187     100O��u��SQ�rzV���\;ȗ��j����d�x�&F��  �b��;����%��m�)+'$r/���è	�q�(aG�H��wi�ԳU��B�z[�Q��5:����ǚ�י%�E�]�E�b��K�^�I��w���U�������1�Y��3��Ylū���
o.���}ޘ�F��w���f��B�1�yE�M�&�����`����iS���~zNpt��b���Cʷ�Y:�!�{���?j�_7����V