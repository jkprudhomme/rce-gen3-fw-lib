XlxV64EB    1054     6c0�ʪҙ��V���Pҍ9�2٫8��A����Vn.ib[w.��mÞ�|��e��^�!����l2u2�%�D�B��&����W>V����7m����贝i�c*���o6:ŦB�	j��������Xαt�b���p@��^ț94���~�=�@�&^�`M>�c��2����iN�Y�����7�REu�Q4���!�8t0%�$��2PZ#>���������;|����0�����%��>V���sNF?D�*���������S��V���FI�%ꏪ��9��kd �!��f�^$3���4�� ��b�i���T������;�T~��N��]Ff��W�=l��R��?�<	#����!�9���9BC`���Ӓ���3zZ�gZHyJ6�L*|y�ڏӎ��Yr:��^$*�mD)�M^����N�F:�� �%�^k�����L��p�����T�����-Vs��N=)��(j-�U��j	%�����p���qV|0ϡ�S�:�0�}��o�V`�&Z�&|�F��ඥ\F�~Бw�fe�V�w%$�|_�BNf];����z�&�K�l�j{�D�lG�P�)��?����:�7<� ����!O���� X=8^��P�X���d"�,GՆ3�aiG{_&ٟ(��/]��o�A�Q�+|��|���W��gꨏss��G�IC{��ұ4��bm-��C`bk��d�M��<��كW�d��ʹ�l��H�����z�1�G05��L)c����<�Ư�S�m��Lz�օ�q.�$
�^va��)I��Y�8 �s���4Wo�(�cc H�6��<��E�zѫJgN<�ƺ��I�t���s0�s!/Q!�9{E+<[� O뗶�=�ӳd���F�!`=
�N����pR@����eW͵b+tV]셡��4KO����-D�Q^�s�W2'��M�<ܔFD
 oM��;�_�c{r�*G��l5��N;B�����q�N�)K�i l7��+m�y��Vh�;fЖY�P*����բ���ռG�M�HM�=�U���}eDp�2
^n��!.�q�|��큿�*5�<����SK�oh\1اaj�	|7�a峔�� u����b�I_�g�3=��ة�^�gY�>���J�}��3!�wͤ�ߐ_����g%�Y�>��m�����ʦfF9���Cۦ:�%C�"7��\�I�s�1Î7{��e�� ȕ>Խ��Ow���Ʒa�qm��Q�K0�m�#�L%���^nN���TXߺy���y�M,V�`p�������z��ԧu��6��>�	�fə\��+?Mb>�9Qĳ��8׹Է�b��A5�R�"�m��"Ts��Ƈl�HV�i.�^�Ow�=�Kd�h$6M޶���#���PY���� ��D�ݖ$P��X�5,�����	�4ĺ
"NQx��|����-�W ���k�Ќx�x"s45ȴ����ou	�#�R	0�T-�m|�+)W�o�\YHMiu���j^oܽE�5O�E2�W ����A�8脠73d玆dc�O���
�Ss��o������֧7�@.O���́�^�{��m��,�L��� 6�^y�4�L�_Z�o~�P8�H@�*Ժ�����>��*�4l�0�k��Z�Aɱ�].�QW��}[6I���o��(�9��шV�6��.�Na�go��~87 _���/�N