XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     170��Y��K_͝G�r9��cxRM*�+�)�IJ!���j����x���NA$B`�A�Y�Q;M�"kJ�f7���i�gd�6�m�ȃ�6;t��pJz�����V3���.��T��d�b�z��-�� W4�P�������Y>M5�	t�^v��Y��)�k������sĿ�d������=��hX��-w���ҫ�a����P{=���}O�����æFy���&����H��:t_��=�*eE5|�]�1�3)���m��n��̣r������`�w*����ul�����x	��Ć���t���	���;�!%)�qDI��<ݒ�{����M���q���8?�����KV���(j��f<i���mXlxV61EB     400      c0�+���8�QP,'
J���UR�ӡ�|l�X�Z�Ѯ$d��_�F4[�5Lk�.�Y��U7�#�����6<Z�l#�c ܆$�pl�� �OV��C��3��NZ!��;0��,�)⩍Dfh.s����<+��%��ౄ���
��?���D�&�_-`��	i�F&��5R1p��099hXlxV61EB     400      d0Ȭ�Qu���1Ĉ�s�Ȫ0k����76����=5}�t�9E����ޡ|+���[]@j"3��a&��"�0͔���#�K�� �k?Æs
�)5ԀV�ˑ=@�ю'?�d�s�#�\���;˃/+a��I�!6�u�'�dB`��D^�<�	�x���"�sᶠV)|�$h{�+��t���n�U����5dp�ܜ(��<�ʁ>Y��XlxV61EB     400      90�<Y��6���D��AD7u�Y���d��ؚٻߔ�d��%�ǂzH7�f(u���Y q/��g�~��\�⥽����M�:���%΢1E7�YG�IK\�����n����y���;�>��\�3�����>u�}XlxV61EB     400      b0FNmQ ��"6���@�G�os.��,�8�g����	���,�Xy�F���v/d�w�+���9�{o#���Z�0��,��0&������ ���Ja�&b�"��)�����ݭ!��g��[5��#��H�8��x��X2�(�S�}��z1e�{o�� �:�aC����:�rA�XlxV61EB     400      90^���ab��R�d�U��M�|EY��D�܂�<��g�'|�&��0� �+�� |V�q�r��ߪ���}�J9�����Xc�:���R�ba�x�#����l�[��_[��x��^��s#�AB7���q�����Ay�H�F����o��XlxV61EB     400      a0���J���P��{Qܯ������Ә�ʧ)H�O<1�x4W����sG�2��L��&��� t�z� (hz�kPYL��L�����O�'v�ʚ��_������t��Jlmf�o�7����M��y��|����5l�v���|��B��"�E��0>��XlxV61EB     400     110+������l��ӽ!�s��RL����| ���p
�����'s�'�=���d���\l�f8�����_�Z��4Z�@�� L}�'��RH�ɬϫ�fGK��+([���.J�m�/1$[k�T,K����q���brW������)���0�vB�a��b?�b$��dRtR�uO�Li�l���	��!��"^�~���������FH5ZpN��5on���)�.�M�eR������>��!��������T�G:9�Um�� �滞��Hg�0��,���XlxV61EB     400      e04zN����՞㯄�\~M��Y13�[Ec�gcvi�����zNSA
5�50�T�6�-7oed}j���Pգ�C��Z;�y�)���NgG$ˀq���<��x���C ���+bZ»(1bn��v�ò�ϕ5;�����d�T�Kjh�[�	~z#�,w#��D>�eݐJ���51�tՌ�v[��"W���$!��V��@jT~:��O^S�Ry�&��`W�4�P�XlxV61EB     400      f0�I�k�;q�PXh�N��*%k�����{��X�` �v*x�Pן��@��\K>�3[)ߗ_� ��
o���t����K������_��F<�� �}�oN@Tڇ
��|@�!��vO?sf��z i��O�r;�D�ќ��<ҳFH���Lhc���dC[l�/-��h��^s�m���@��-
����D�!����~(݀�d��L���:��TN�ʋ�B��#�~�0�u�&����w*O�XlxV61EB     400      e0`���V�4��?4�deQ��/V���4�-��
@��/
���+�H�p�1��Hu�a(�TkG����`:ee+v�"�j*��xX�5�p�	���0�P�a�E�aL��D�:*L��6adaٟ�����!��CH�����r�y������p?èK�� p��ڎs�4�����@�=��D�b$�7�v���VԹM#�G[��<�K	8�:�P�-�	�?%�ΚXlxV61EB     400      e0x���0��j�3?
šW�x������U��6�%��F7���Z|ϔ0h�O:�-���i:&+m%�GF6�Z3n�/�`��q�`��������������g;[�=�t��#~N�1�;	�Ƥ�"Y)R�� �|����\Gխ��vZ�?i=��4ƽ���S)���E��UA�/\(j/Ze���Pf�����P� �X��َ�GJm[܂�+U�4 �bD�`XlxV61EB     400      e0Q?!�9��`�Hl���@x�աU_l� �"m(�l?Ϟ��ʑA/ٮ :E��
���)��~�<�޵��Nl��ai����t[�e��d<�����궛�Qz�?����-6MѺv%+4�K�[���Y���0�����e�A溘5q��)��L���-�%�����U��p��7�3}s[@Qf�	g��*W�=�s��j��[���N[p~�c�j���>�q褟XlxV61EB     400      e0G�awn�'���.fEr��JAL�'}p�$� $�'�K#�;1�[�A�پ�o4�:ˇpȉ�� u$ ��/�ǵ��S���&�;�X([�HҸ��a��w�~GjqI�����ec�/�Ā��=g���'�������/#�;�P:�V����;�x��y�tDq^	-���Q�5џ�_9t�ӄ��ş�l��-|bA��M\�jNz�\�ޝ�ꨏrAXlxV61EB     400      e0HnQ���{6b����]�C��^K�}�x��8D�+�+�K���L���z�d.�3>,�tW8x"�y
C�2�A;�AF|x|p��A���*�o�vg�fѓ-A;�C����_NQ�O�2�܁;�G�qΉߤ~�v�^v>�.��K8N��U�~ΐ6)ɔ�����ϒ�78>�$q�r�R��.__�(���FQ.NR�����zl`�Ҥl���~��XlxV61EB     400      d0
�VX��pU')0�;2�VW3�?A�]?;2s��������.�`��9�r���0������AX���z�c�q�	v�j��\�c�EV�#?'9H��؀xZ���]�&�"��Հ�m���1 �\�,��ӧ�o'��}�LC�̰+���7`'2��0�=��t�S��l5fz8K����E�,�fP��.u/��v��t�Db�&iXlxV61EB     400     130�:F�����j�y��kidp��tG�����,�Þ���o��2�";��ڇ��:l���E�'��A
s��Y����U�;��;������R:����4(T:G�ޔ24o���:}�k�3:wB�t2����H��3gZ��?m�,�^�i��:^X�準ʀ�j�T~R_�ޒ�U#�ȀG�2r�r}�)i�n��1i���qc�/�l
w�>;�|0����2�n����έ�@�HӋ3}�����r�D�Z>m���,��gf�N���p�=��o@�Z8��H�.2/���e���@hXlxV61EB     400     120��{aE�������ۨ!�Å.�r� >hE`d07�G�ؾ�o�3�ؑYO�.��Ó{�+ӞF�#1����T���K��x|��K�4E�"w"���Ed��Ƴ*��%��H-N��퍴��ׄ�6K��)��-����	��wց�C	��^H�*��������p�!��Vvaw�d�P	�o�x�K�5����
_�|�p|$� O~T��>���D�C&A�4h=��h!bf�3���9vM#Y?��'��J�� Uh��5\%Sb�ᡴp(EK�N�^G�KXlxV61EB     400     140�tST�����X��YV۱8���_�.�� ��|�"aE�#ln��JsA��,���� r��N�Z��#EX�l��E��aT�"$�O��?�Y��o;��?H#�6����]y6����)��.���M[����>L)��v��7u7�J\�\��4���2�(��k�!傋�%�O};%�δe�} :Q���V��f"E9�����x���:�g9�{9����J�YV}#��Xč�u�Y��ɵ��g3�/��JIsz~������}��\\T�/�p�0���DbE��2���� �?@8B�^	�t�:�t�D�����=[XBx1XlxV61EB     400      d0�D㼎)�[�)�VUv���ks/�w��U�4��v5�2sm��+]�j�ۅ NJ�m��ĺ�AFe���`���dd#�S���Ý����p�!�1�{�M��h���(}|m8g���{����^��}>q�2��ǵ�g�'��Y�>_��k��p�l�^દ�Jw�m�� �{�����(�]^��wa��
�k�Z�s�rY���:(]�O�XlxV61EB     400      d0SO�G+��,)��P�����]H��lS �Ԑ[�T9^������0�4���/4vȀ�ł���uU�U�7gQ���u�\�,�o�«<0���BtPr���9��DD�"ر2_�0����ACא0����`���H�������ǻJ-�=��S-�]�V�d�-���=w�j4
!rߢA��=���&��ZL��������XlxV61EB     400     100�C�L�)�Rop�?p$I�o4\�H�l���3m[A�=�-,$:�**1MI��ZL���9��_��d�B�
N�C��<*�bM�R�E�+Z&���cj��q��o�[I�H^��������W���e�m�Ce��n��ڀ�ȟ�l-�����I*ސ`��%%&өn����$!�6���~K���/0"e$r� sn�S^��F`V�����N�4Q^�T��M�'�ѬS�>6H��'�c�Y `\'M�PXlxV61EB     400      c0:T%`�d��(�[L�J�8��[����t��q&��
?�PM�hH��M�	��h9 ����J�I�ò\<Z�#Gs��-�
��	�n9:�P(O�����^�w^�_��^����>&���p�l=xz]F�5������Dh���<mE��SԪ5k���7�A���Z��M�:=�b���a�0|XlxV61EB     400      c0� ��Qʀh]��*b��K(Uɡ|9�ݏ��U���b�py�����^fh[9��Uh�0Ѳ�&@(�~Vf@{'���C�~W��U�^���[n�K�
ǓW��%���!{J�m{	�n$F���9
x�p���l�A��җ��R�;�ؿ��c�Zi��Ł\%0Շ�� ���������1P�Dp��[H۲�GnXlxV61EB     19c      90��X����2�����%Fâ�}���wVV�Ee������W���ǉ�4!��(��K������Ы~�N�ԩ'�����gz���� �����)!�t+�K�i��Q�&E�p���K6�����8"!��6d9��}��;�,