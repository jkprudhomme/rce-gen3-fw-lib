-------------------------------------------------------------------------------
--
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : zynq_xaui_gt_wrapper_tx_sync_manual.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\ 
--
--
--  Module  zynq_xaui_gt_wrapper_tx_sync_manual
--  Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2011 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 

 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--***********************************Entity Declaration*******************************
entity zynq_xaui_gt_wrapper_tx_sync_manual is
   generic
   ( NUM_SLAVES	: integer := 10 	--Should be non-zero
   );
   port
   (
       START			        : in  std_logic;        
       PHASE_ALIGN_COMPLETE             : out std_logic;       -- Indicates Phase Alignment complete on all lanes
 
       --Master Signals
       M_GT_TXUSRCLK   	    	        : in  std_logic;
       M_GT_TXRESETDONE		        : in  std_logic;

       M_GT_TXDLYSRESET		        : out std_logic;
       M_GT_TXDLYSRESETDONE		: in  std_logic;
       M_GT_TXPHINIT		        : out std_logic;
       M_GT_TXPHINITDONE		: in  std_logic;
       M_GT_TXDLYEN		        : out std_logic;
       M_GT_TXPHALIGN                   : out std_logic;
       M_GT_TXPHALIGNDONE               : in  std_logic;

       --Slave Signals
       S_GT_TXDLYSRESET		        : out std_logic_vector (NUM_SLAVES-1 downto 0);
       S_GT_TXDLYSRESETDONE		: in  std_logic_vector (NUM_SLAVES-1 downto 0);
       S_GT_TXPHINIT		        : out std_logic_vector (NUM_SLAVES-1 downto 0);
       S_GT_TXPHINITDONE		: in  std_logic_vector (NUM_SLAVES-1 downto 0);
       S_GT_TXPHALIGN              	: out std_logic_vector (NUM_SLAVES-1 downto 0);
       S_GT_TXPHALIGNDONE           	: in  std_logic_vector (NUM_SLAVES-1 downto 0)
   );

end zynq_xaui_gt_wrapper_tx_sync_manual;



architecture RTL of  zynq_xaui_gt_wrapper_tx_sync_manual is

--***************************Parameter Declarations*****************************

    constant DLY : time := 1 ns;

    constant TIMEOUT_VAL : std_logic_vector(19 downto 0) := X"186A0";  -- 100K CLK cycles 

    type state_type is 
                       (INIT, SRESET, MASTER_INIT, 
                        MASTER_PHASE_ALIGN, MASTER_DELAY_ALIGN,
                        SLAVE_INIT, SLAVE_PHASE_ALIGN,
                        MASTER_FINAL);

                        


--************************** Register Declarations ****************************
    
     signal    present_state, next_state	: state_type;
     signal    all_lanes_dlysreset_done         : std_logic;
     signal    all_slaves_phinit_done           : std_logic;
     signal    all_slaves_phalign_done          : std_logic;
     signal    m_gt_txdlysresetdone_r           : std_logic;
     signal    m_gt_txphaligndone_r             : std_logic;
     signal    m_gt_txphaligndone_det           : std_logic;
     signal    m_gt_txphinitdone_r              : std_logic;
     signal    m_gt_txphinitdone_det            : std_logic;
     signal    m_gt_txphaligndone_2r            : std_logic;
     signal    m_gt_txphinitdone_2r             : std_logic;
     signal    s_gt_txdlysresetdone_r           : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphaligndone_r             : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphinitdone_r              : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphaligndone_2r            : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphinitdone_2r             : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    m_gt_txdlysresetdone_det         : std_logic;
     signal    m_gt_txdlysresetdone_det_r       : std_logic;
     signal    s_gt_txdlysresetdone_det         : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txdlysresetdone_det_r       : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphinitdone_det            : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphinitdone_det_r          : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphaligndone_det           : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    s_gt_txphaligndone_det_r         : std_logic_vector (NUM_SLAVES-1 downto 0);
     signal    phalign_lost                     : std_logic;
     signal    done                             : std_logic;
     signal    done_d                           : std_logic;
     signal    timeout                          : std_logic;
     signal    timeout_match_d                  : std_logic;
     signal    timeout_match                    : std_logic;
     signal    timeout_cntr                     : std_logic_vector(19 downto 0);
     signal    st_chng_d                        : std_logic;
     signal    st_chng                          : std_logic;
     signal    all_lanes_phaligned              : std_logic;
     signal    all_lanes_phaligned_r            : std_logic;

     function and_reduce(arg: std_logic_vector) return std_logic is
	    variable result: std_logic;
     begin
	    result := '1';
	    for i in arg'range loop
	        result := result and arg(i);
	    end loop;
        return result;
     end;
begin
--************************** Beginning of Code ********************************


    --__________________ State Assignment______________________________________

    process (M_GT_TXUSRCLK, M_GT_TXRESETDONE)
    begin
       if(M_GT_TXRESETDONE = '0') then
          present_state   <=   INIT    after DLY;
       
       elsif (M_GT_TXUSRCLK'event and M_GT_TXUSRCLK = '1') then
          present_state   <=   next_state    after DLY;

       end if;
    end process;


    --__________________Next State Generation______________________________________

    process (present_state, START, all_lanes_dlysreset_done, m_gt_txphinitdone_det, 
             m_gt_txphaligndone_det, timeout,
             all_slaves_phinit_done, all_slaves_phalign_done, phalign_lost )
    begin
       case present_state is
       
       when INIT =>
       --START indicates DRP write to X06F is complete and Phase Alignment can begin

            if (START = '1') then
               next_state   <=   SRESET;
               st_chng_d    <=   '1';
            else 
               next_state   <=   INIT;
               st_chng_d    <=   '0';
            end if;
   
       when SRESET =>
       -- Assert TXDLYSRESET for all lanes
       -- Deassert TXDLYSRESET for the lane whose TXDLYSRESETDONE is asserted 
       -- Wait till TXDLYSRESETDONE for all lanes is asserted

            if (all_lanes_dlysreset_done = '1') then
               next_state   <=   MASTER_INIT;
               st_chng_d    <=   '1';
            elsif (timeout = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   SRESET;
               st_chng_d    <=   '0';
            end if;
  
       when MASTER_INIT =>
       -- Assert TXPHINIT on Master
       -- Deassert TXPHINIT on the rising edge of TXPHINITDONE 
            if(m_gt_txphinitdone_det = '1') then
               next_state   <=   MASTER_PHASE_ALIGN;
               st_chng_d    <=   '1';
            elsif (timeout = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   MASTER_INIT;
               st_chng_d    <=   '0';
            end if;

       when MASTER_PHASE_ALIGN =>
       -- Assert TXPHALIGN on Master
       -- Deassert TXPHALIGN on the rising edge of TXPHALIGNDONE 
            if(m_gt_txphaligndone_det = '1') then
               next_state   <=   MASTER_DELAY_ALIGN;
               st_chng_d    <=   '1';
            elsif (timeout = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   MASTER_PHASE_ALIGN;
               st_chng_d    <=   '0';
            end if;

       when MASTER_DELAY_ALIGN =>
       -- Assert TXDLYEN on Master
       -- Deassert TXDLYEN on the rising edge of TXPHALIGNDONE 
            if(m_gt_txphaligndone_det = '1') then
               next_state   <=   SLAVE_INIT;
               st_chng_d    <=   '1';
            elsif (timeout = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   MASTER_DELAY_ALIGN;
               st_chng_d    <=   '0';
            end if;

       when SLAVE_INIT =>
       -- Assert TXPHINIT for all slaves
       -- Deassert TXPHINIT for the lane whose TXPHINITDONE is asserted 
       -- Wait till TXPHINITDONE for all slaves is asserted
            if (all_slaves_phinit_done = '1') then
               next_state   <=   SLAVE_PHASE_ALIGN;
               st_chng_d    <=   '1';
            elsif (timeout = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   SLAVE_INIT;
               st_chng_d    <=   '0';
            end if;

       when SLAVE_PHASE_ALIGN =>
       -- Assert TXPHALIGN for all slaves
       -- Deassert TXPHALIGN for the lane whose TXPHALIGNDONE is asserted 
       -- Wait till TXPHALIGNDONE for all slaves is asserted
            if (all_slaves_phalign_done = '1') then
               next_state   <=   MASTER_FINAL;
               st_chng_d    <=   '1';
            elsif (timeout = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   SLAVE_PHASE_ALIGN;
               st_chng_d    <=   '0';
            end if;

       when MASTER_FINAL =>
       -- Assert TXDLYEN on Master
       -- Wait for rising edge of TXPHALIGNDONE on Master
       -- If TXPHALIGNDONE of any lane is deasserted go back to INIT
            if (phalign_lost = '1') then
               next_state   <=   INIT;
               st_chng_d    <=   '1';
            else 
               next_state   <=   MASTER_FINAL;
               st_chng_d    <=   '0';
            end if;

       when OTHERS =>
               next_state   <= INIT;
               st_chng_d    <=   '1';

       end case;
    end process;


    --__________________Output Generation______________________________________

    process (M_GT_TXUSRCLK)
    begin
       if (M_GT_TXUSRCLK'event and M_GT_TXUSRCLK = '1') then
       case present_state is

       when INIT =>
               M_GT_TXDLYSRESET       <=   '0'    after DLY;
               M_GT_TXPHINIT          <=   '0'    after DLY;
               M_GT_TXPHALIGN         <=   '0'    after DLY;
               M_GT_TXDLYEN           <=   '0'    after DLY;
               PHASE_ALIGN_COMPLETE   <=   '0'    after DLY;

               for i in 0 to NUM_SLAVES-1 loop
                 S_GT_TXDLYSRESET(i)       <=   '0'    after DLY;
                 S_GT_TXPHINIT(i)          <=   '0'    after DLY;
                 S_GT_TXPHALIGN(i)         <=   '0'    after DLY;
               end loop;
        
       when SRESET =>
       -- Assert TXDLYSRESET for all lanes
       -- Deassert TXDLYSRESET for the lane whose TXDLYSRESETDONE is asserted 
            if(m_gt_txdlysresetdone_det = '1') then
               M_GT_TXDLYSRESET   <=   '0'    after DLY;
            else
               M_GT_TXDLYSRESET   <=   '1'    after DLY;
            end if;

            for i in 0 to NUM_SLAVES-1 loop
               if(s_gt_txdlysresetdone_det(i) = '1') then
                 S_GT_TXDLYSRESET(i)   <=   '0'    after DLY;
               else
                 S_GT_TXDLYSRESET(i)   <=   '1'    after DLY;
               end if;
             end loop;

  
       when MASTER_INIT =>
       -- Assert TXPHINIT on Master
       -- Deassert TXPHINIT on the rising edge of TXPHINITDONE 
            if(m_gt_txphinitdone_det = '1') then
               M_GT_TXPHINIT   <=   '0'    after DLY;
            else
               M_GT_TXPHINIT   <=   '1'    after DLY;
            end if;
 
       when MASTER_PHASE_ALIGN =>
       -- Assert TXPHALIGN on Master
       -- Deassert TXPHALIGN on the rising edge of TXPHALIGNDONE 
            if(m_gt_txphaligndone_det = '1') then
               M_GT_TXPHALIGN   <=   '0'    after DLY;
            else
               M_GT_TXPHALIGN   <=   '1'    after DLY;
            end if;
 
       when MASTER_DELAY_ALIGN =>
       -- Assert TXDLYEN on Master
       -- Deassert TXDLYEN on the rising edge of TXPHALIGNDONE 
            if(m_gt_txphaligndone_det = '1') then
               M_GT_TXDLYEN   <=   '0'    after DLY;
            else
               M_GT_TXDLYEN   <=   '1'    after DLY;
            end if;
 
       when SLAVE_INIT =>
       -- Assert TXPHINIT for all slaves
       -- Deassert TXPHINIT for the lane whose TXPHINITDONE is asserted 
            for i in 0 to NUM_SLAVES-1 loop
            if(s_gt_txphinitdone_det(i) = '1') then
               S_GT_TXPHINIT(i)   <=   '0'    after DLY;
            else
               S_GT_TXPHINIT(i)   <=   '1'    after DLY;
            end if;
            end loop;
    
       when SLAVE_PHASE_ALIGN =>
       -- Assert TXPHALIGN for all slaves
       -- Deassert TXPHALIGN for the lane whose TXPHALIGNDONE is asserted 
            for i in 0 to NUM_SLAVES-1 loop
            if(s_gt_txphaligndone_det(i) = '1') then
               S_GT_TXPHALIGN(i)   <=   '0'    after DLY;
            else
               S_GT_TXPHALIGN(i)   <=   '1'    after DLY;
            end if;
            end loop;
   
       when MASTER_FINAL =>
       -- Assert TXDLYEN on Master
               M_GT_TXDLYEN          <=   '1'       after DLY;
               PHASE_ALIGN_COMPLETE  <=    all_lanes_phaligned   after DLY;

       when OTHERS =>
               M_GT_TXDLYSRESET       <=   '0'    after DLY;
               M_GT_TXPHINIT          <=   '0'    after DLY;
               M_GT_TXPHALIGN         <=   '0'    after DLY;
               M_GT_TXDLYEN           <=   '0'    after DLY;
               PHASE_ALIGN_COMPLETE   <=   '0'    after DLY;

               for i in 0 to NUM_SLAVES-1 loop
                 S_GT_TXDLYSRESET(i)       <=   '0'    after DLY;
                 S_GT_TXPHINIT(i)          <=   '0'    after DLY;
                 S_GT_TXPHALIGN(i)         <=   '0'    after DLY;
               end loop;

       end case;
       end if;
    end process;


    --__________________Internal Signal Assignment___________________________________


    -- done indicates that rising edge of TXPHALIGNDONE in MASTER_FINAL state

    done_d  <= '0' when (present_state = INIT) else
               '1' when (present_state = MASTER_FINAL and m_gt_txphaligndone_2r = '0' and m_gt_txphaligndone_r = '1') else
                done ;


    -- Timeout Logic for each state
    timeout_match_d   <=  '1' when (timeout_cntr >= TIMEOUT_VAL)           else '0';
    timeout           <=  '1' when (timeout_match = '1' and st_chng = '0') else '0';

    process (M_GT_TXUSRCLK)
    begin
       if (M_GT_TXUSRCLK'event and M_GT_TXUSRCLK = '1') then
          if(st_chng = '1' or timeout_match = '1' or present_state = INIT) then
             timeout_cntr   <=  (others => '0')    after DLY;
          else
             timeout_cntr   <= STD_LOGIC_VECTOR(UNSIGNED(timeout_cntr) + 1)    after DLY;
          end if;
       end if;
    end process;

    
    -- Logic to detect the rising edge/ assertion of various *DONE* signals
    process (M_GT_TXUSRCLK)
    begin
       if (M_GT_TXUSRCLK'event and M_GT_TXUSRCLK = '1') then
           m_gt_txdlysresetdone_r       <=   M_GT_TXDLYSRESETDONE        after DLY;
           m_gt_txphaligndone_r         <=   M_GT_TXPHALIGNDONE          after DLY;
           m_gt_txphinitdone_r          <=   M_GT_TXPHINITDONE           after DLY;
           m_gt_txphaligndone_2r        <=   m_gt_txphaligndone_r        after DLY;
           m_gt_txphinitdone_2r         <=   m_gt_txphinitdone_r         after DLY;
           m_gt_txdlysresetdone_det_r   <=   m_gt_txdlysresetdone_det    after DLY;
           done                         <=   done_d                      after DLY;
           st_chng                      <=   st_chng_d                   after DLY;
           timeout_match                <=   timeout_match_d             after DLY;
           all_lanes_phaligned_r        <=   all_lanes_phaligned         after DLY;
       end if;
    end process;

    process (M_GT_TXUSRCLK)
    begin
       if (M_GT_TXUSRCLK'event and M_GT_TXUSRCLK = '1') then
           for i in 0 to NUM_SLAVES-1 loop
               s_gt_txdlysresetdone_r(i)       <=   S_GT_TXDLYSRESETDONE(i)        after DLY;
               s_gt_txphinitdone_r(i)          <=   S_GT_TXPHINITDONE(i)           after DLY;
               s_gt_txphaligndone_r(i)         <=   S_GT_TXPHALIGNDONE(i)          after DLY;
               s_gt_txphinitdone_2r(i)         <=   s_gt_txphinitdone_r(i)         after DLY;
               s_gt_txphaligndone_2r(i)        <=   s_gt_txphaligndone_r(i)        after DLY;
               s_gt_txdlysresetdone_det_r(i)   <=   s_gt_txdlysresetdone_det(i)    after DLY;
               s_gt_txphinitdone_det_r(i)      <=   s_gt_txphinitdone_det(i)       after DLY;
               s_gt_txphaligndone_det_r(i)     <=   s_gt_txphaligndone_det(i)      after DLY;
           end loop;

       end if;
    end process;


    m_gt_txdlysresetdone_det <=   '0' when (st_chng = '1') else
                                  '1' when (present_state = SRESET and m_gt_txdlysresetdone_r = '1') else 
                                   m_gt_txdlysresetdone_det_r;

    m_gt_txphinitdone_det    <=   '1' when (present_state = MASTER_INIT and m_gt_txphinitdone_2r = '0'and m_gt_txphinitdone_r = '1') else '0'; 

    m_gt_txphaligndone_det    <=   
      '1' when ((present_state = MASTER_PHASE_ALIGN or present_state = MASTER_DELAY_ALIGN )and m_gt_txphaligndone_2r = '0'and m_gt_txphaligndone_r = '1') else  '0';



    process (present_state,s_gt_txdlysresetdone_r,  s_gt_txphinitdone_r,  s_gt_txphinitdone_2r,
             s_gt_txphaligndone_r, s_gt_txphaligndone_2r, s_gt_txdlysresetdone_det_r,
             s_gt_txphinitdone_det_r, s_gt_txphaligndone_det_r)
    begin
           for i in 0 to NUM_SLAVES-1 loop
               if ( present_state = SRESET ) then
                  if(s_gt_txdlysresetdone_r(i) = '1') then
                     s_gt_txdlysresetdone_det(i)    <=   '1';
                  else
                     s_gt_txdlysresetdone_det(i)    <=   s_gt_txdlysresetdone_det_r(i);
                  end if;
               else
                  s_gt_txdlysresetdone_det(i)    <=   '0';
               end if;

               if ( present_state = SLAVE_INIT ) then
                  if(s_gt_txphinitdone_2r(i) = '0' and s_gt_txphinitdone_r(i) = '1') then
                     s_gt_txphinitdone_det(i)    <=   '1';
                  else
                     s_gt_txphinitdone_det(i)    <=   s_gt_txphinitdone_det_r(i);
                  end if;
               else
                  s_gt_txphinitdone_det(i)    <=   '0';
               end if;

               if ( present_state = SLAVE_PHASE_ALIGN ) then
                  if(s_gt_txphaligndone_2r(i) = '0' and s_gt_txphaligndone_r(i) = '1') then
                     s_gt_txphaligndone_det(i)    <=   '1';
                  else
                     s_gt_txphaligndone_det(i)    <=   s_gt_txphaligndone_det_r(i);
                  end if;
               else
                  s_gt_txphaligndone_det(i)    <=   '0';
               end if;


           end loop;

    end process;
      
       all_lanes_dlysreset_done  <=  and_reduce(s_gt_txdlysresetdone_det) and m_gt_txdlysresetdone_det;
       all_slaves_phinit_done    <=  and_reduce(s_gt_txphinitdone_det);
       all_slaves_phalign_done   <=  and_reduce(s_gt_txphaligndone_det);

       all_lanes_phaligned  <=   and_reduce(s_gt_txphaligndone_r) and m_gt_txphaligndone_r and done_d;

       phalign_lost  <=  '1' when (all_lanes_phaligned = '0' and all_lanes_phaligned_r = '1') else '0';

end RTL;
