XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     140���<&45�܆��>/�Y�.5*���pNlń�/
�%�j#]Z~]���)�tI~�y'e+�K��mͭ��$P��xN:v"�R��d>�-���GI�[a��p�F	tpD��|<��		�y��R+�N(��z���=;��#�7ʯ�G��-��S��Q�ξ7K��b��b(�Z
��
�/\D�t"��K2~�K�b�����ړ#�x4�V�0��$����)�)J(���:ɒ��kVPD�6o�J��
r
��"��T�HS��O=C`mӭ�xK)!%�䎋~�.��ʨ����@��G���&8o��|@XlxV61EB     400     1a0qOU()p8�e3���G���	�
���� f� �b:Z�s����6�Z��t�8;�
^GW�۫��Ho�r�U���I�U��IO8͠�2�E3`���1Q�H�w+�J|ê�|��=�f��3_q[��\�lL��=ǹ�W���	!��LƌF�n���� !%��J5�6��>^,>~ob
�kK`͠�~��V��q�'N�����iH�%V��8�e�⮍ZL��X~���U�+�S�^�(�,��JA`���χ�P�Wsg���-��nײ�JaiS����oC�&J3h{�
ZH���.�L@5�@�7ċ+�("=ةӯ�]���Z���6?:���d��S�����ZG ��L��
\w�� ��ܵ8��$e��]������T��a�y_;͸T`�ϼ"0ܿX�hXlxV61EB     400     180�����%�c��1���os7T(�r���5N\�V8�2oS���*q򾅣	2�w_�v&�Q<�V���jF�cž�S8��6�-�~�Bꠀ��DM���[�ǃ���@�J��Q�R�D�{[.%���^9Ѐ�/,� ����f��֤m�u �P�Z���"L����E�/ 5sU���w��;����r�s���qC��)-/T)���o$屭�/"$�Ƥ�p%�$�.�U�O��`J�g�ql^(���	h�>ϵP�oxǧ3����T�Meװ.	��x�ƽ.F�"^��l������������o@ ��W>�tu�N������1��k�����i��Y	. ;�3���L%�h��
�w����>H��/�7��XlxV61EB     400     130�޹���xC��v<ߎ���p���tFzb���tm���Y�_39������9X�����?��&�P_���!.�yF��4rb��S��lG������ ��s���3���˃��\G��~�A�����S�G�ЮH~9�mЩ^k�(F�X�T1��۵j�7�>�FC�FAKZe��uO,��2A����GR����lՄn�}�x�����A�
S,M+UZŐ��4��kѶ.��L~�ǔic�Gw`/⚑��� 5I��2�W�����8D�p�Α+����rn���-�y��Y
�>��c�c��P�XlxV61EB     400     100�s�֡��Y�	�~&�9���(�ϑ9��o>�,��R�9_���o����ZΠ��Ygna:�>D���(���{7�Aa�hۋ��Rx�G#���p���K�0A`f���s���n�3�o-�QS�XH���r|��&��hVv�/���M`�=m�Z�y6�J3�ٕP�Ϡ/.�2�;B�&ԭ��
��y���R�.TL��zH�)��D��{1�`d�X����D�۠x�`�&v�E�_m/�|k�(����"XlxV61EB     1f7      f0�#���g����bG�S��UiA9��1�D�9�+�����n��ۭ�$�cψ���-#"��%�F�ĥY-�7�q�h8)�w�.w ➑�i����q�:)�΍J�B���I�a�az?��K��R��ڤ��uV���`L34��M'������Z}��bRw��1ي����o~��zEO�����
>׼�����)	O�(d�w�p+<��e��:~H�~��f�,8���h�