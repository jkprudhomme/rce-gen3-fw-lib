XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180���G
Ø"-�Y��	�lo�Nʈ LM|R� w%=~V��-��y1F���~�����#@"Q��U\J.���Ow�����É���ާM���Y��[ŵ����"e�M1j⪍���7�=�?>o��0������&}Y\$&�K�1�o��m�{+�X�e(��`��Yp�{K~��J����)���Q~a�v{Ëo����C?�݋zl�E3�>�޶����,��z���1��G�Q��]����"y�9?���s��TA���ӋE���L�`U�lJ+L69����reB㨀��u�1i9f�L�|�뺢��^)2���Z�g��2Y[ �P�;�~�g��^{_�^S�zS����S!s�p�X���S��@�w�u^&+�B��g	XlxV61EB     400      e0�
�l�+��E�����8 )��Ѿ��WА��|�`���=��E��*�����Qn��;`ڢ�GY6C��,��(�2��W\���&��B��ç�{�T�dF��ۄ+��Ұ�����"1�E٨��E�f0�<��}S:QI0`j��9�����i�)c5�D��9�Ɋ���p����^�@�.���8�g��G�_�~��z�\%��g9Z��� 0�?XlxV61EB     400     140,aMP@o������Wɫ%;~,ȼf��H���끗n�3�sg��5�U�|��S�q�O������,� X3	�_��%m�Y��e��,�B���j�W����ߋX��~�(��fR�!�l�wx�!Ռ��^���F<��{��F�MnE%��� >Y��ؒ�0�B�D�6�de1Ņ�
D8F@���!L�;7��rc	�ĦR��X�K��dIü��m�����8�N���l}o�k$?��Lĩ�UU�5)��ĳ��戫P�Q���A� R���Ƅ���})�������e�x��R9��AJT�.Pps#XlxV61EB     400     190�Vx��??����%5�����qD	�ވ�8@���ݛb�h�r��D� [���},, *}�h��C��`�����W�[v��U.�bB�TΉ{�/����"��>͞��VSrģ�nK�=ja-��.���
	n5�~�԰<fV������ q��@,�����zΪ���aK�=s��6O����+�.��Dz.�'`�83����bJQ�J>B뤭-%��b��m�������ާ�t2{����I@M�x�= b�Zd�U� ^��'4������oو��i�0gL�8�ǦF��Gہ!��)Pv�aVՀ�'J�an�e/���f����Dm�=��	)�Ʋ?��
U�_��|3�壉��BBi)a����С
.=���v&xnW�ʏ�[5y7eS��XlxV61EB     400     100��a�1�����X��4��i"F�|(�>�8b�������(%B����]"�;��[8s�� �^���㯿=s"�a$��¦�F�p'����@b��9冹?	E)�Ś����e[�kIGE�^b��c�He.��p�x�x<���@�v�)2�Dh̗��Y"�_ۃ=>jk���3n�ל�Mv1ö���+A4Cꞩ<*� R��$᷅��p��g`�ki?@�z��3^�90J�c�z��ģ�]g��XlxV61EB     400     110x���[a3�Z	q���������Wktw8��>�a�L����4��� �/�v����L
�i{:�ߴ�n�U��*����+���?�����Z�J�ݐ���M�ľ�C;x�P�]!��[й ac�X(������E� ��|���'����^�0�4��`���[����ҥ��#�/<�-�@[������댿�a]H��B�w�z7���F�Y �1ʠ,�tw��󈁺������V0��i��]{�Z��7k�m�H�r�T��?�V�QXlxV61EB     32f      f0.oihg���z�c4�̻�h�5&��/�r"�'d	�h	����Q�=N��m��O�Z�"��r����-FHm���_B��C�ÿ�����t�����@y�A���/zj��bww'�ppm�!��k6��O�iv���ai��-i��n�j/�F:��'-�V�b����XX�a,����i`��7^s3%��P�XR���m����,c�cp
��yY��Hx�/��b