XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150JviM��	%�ٳ��t(g���:��a������.�~{�17�5�$JG�;�Ho��U�j��eb\�]��}��+�f'|�Z����P���0O@��m�bm��������BIZ���i��9�W�0�p�scȜ�]&��ur
U��.�u���?�
�M��L	9�l�[�91ɻ݅��ן�@Nܬ�I{{0�<��~��@�����{���R���X���4ؘ��AB TS�\�� D���?��G�PA�r^k��Ks�8�(�n����#OPz� bEF���m��W�t��	�t2B�0L���Q4��ܜrK<��,�
E��6�XlxV61EB     400      e0�P��:U�8c�r��)��*�r��U�M�����Q'!�a�{C����+hl�j@��ބ�����X���[�ƿđ,H��g�|�h4��Q�#�8�T�"i`��@�8 a�>݋����w2(�I���vc1k�PX�����,!ǧW�����F�o�����b��)�{��^z(d������~��?���&������L�����`�N��XlxV61EB     329     100�+ �S��и�G��p�^!�]�+��ew�,`}X��}�쟨���#�䌅f���q�z%�~��tPm
Z�GTظ�"a+���f��L��WE�AϮZ��+��8k��$�ql"��jN,���L��(u��GZ�w�㑊�f��ݽ�,[�	�:���FJ �q��\﫰Z�?��8ӝ{g�1��g�KH
_@����?/LB��� ��F�{�6e��� X��)�sG	���>�����@F�v