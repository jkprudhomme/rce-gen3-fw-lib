XlxV64EB    21fb     da0ǣĲ��A������m��}$-�y���A�� �W�o����߹O�@-�'��b!Av6x8��J��P'瀨H"��;�e2�j�i�������r�X=U ����^a����bI� ,�>:O�� F��(iT����S�+>Ddf��K�M�=���?�K���b�\I bb�u�#c�fpqG��A�t���HP��I�,��r ܄�����	}NW�՚�9{� *���bf�)�!&��j����_b�>_P]���̀��5�p����t�Q����2 C��3�ybO�d��7V�X阔A 8�L^T*K�2|�8�����+��=)���&�Y���?Xxd��۵�v��B���U����Y�G��Z<,(avj900@b�M������B�ߎ��4�>��S�2�`���t�&��`T�0���`
���/{R�7�~vi)Dv��Çㄚ@|ǹ�] �+��F��)�i����@j@k��5���vI����c';;�~;��g=tѽ�y����&DU�~�~1_$9|��Bn�Q%���D���J	9�}0z�\.�5��{����˶>ڂ.�x�&�A
�Cw���,p�2��;�!.F�I�#a�b�r��}�ڰ*�%U��Gg���q�ξ�b����
d�����ѥ�	8�'I�j\�O
ʱ}��7��ƀ���b�ǅ�=^���8�]sU �1�:�ku��K�@������z�D�{�T~"����as�{�"�vp���[�z�n)��P�����&��f{(�tM������������u�iy9Ai%��c�0+}B�U��:����!#+S��R�s���p=�Ou�U����`�^��
���0�g���*[�Mr.�kw����p��ٛ�Ю���v��,@��vظ{���-�~`O޳�h����XQ�_�=`y��*W���ғ?��= ��6�)I��4� �}�߲�0;�i/��gc�Й�����qUp%�c�>�g�.w!اc",��'o��>W
L���T&��x�o��aM��l�K@P�C�+��]d0&/.�:�JӦ�w��3���;�s߳�����,��%�5���4�iF�n��T�ͺ���N��,�P�D�|y~�!wBsV�� d+�U�S�n�m���D-��Fg`����/ ��y� �e��A���{�2(�S/�2/e�vF�<�3*�mh��o��P�\�J*a�,��5*�h�|50XD>K#ػV��]�T]y���M������sQb`�6@*��|��fb�~���M�2�Q���BX�,�F��������j	6��AШ��u{�Ν�����|�� I��7*H˨q�� �'���� ��H��̈��ޘD����95n�s��T���Z�HV8�Ĩ����bg��y� w��Z.����lsQ=+�U��~�6���M+����P�A��V�dw�1\k(;�������e�I�:��{>rr6��������dt1��o�>�d9ih����_��8qX,z �*�h�=�)��#�u<�"R�@���t��)j.;n�[�eĀ�nr�ﹹ�߽6�M��w��CE�vFd�<�D;jM�{����m٧���0��U�`�HvX �L�@�?^Pj�:X���7��(��:��v�폦1��w�p{ƅ>Y;z��)�o?�����,�&�b�M�n,�U���fFbQhE�qq���V�1
fȯ�W��]tr{LoAS�^@t1Ǯ�r���#՛5CD��G�eY��:B��
�߮@���n�0�3Z\��]���y��ѧNF���ݨ�r��3���b�����u:):�Oc���qiAAI��@�#R�Y���SG9�V�����`U����0iey���ax����L$�9�/Nb�i�B t�P..�kd��P1��`xˤ�2��2��;�mA�RuND�猑�V�b����� '��U"�R.�6jUӧ�~_�N{~%�i�ۮbl8�@�6Bؚ�bc$��e������25���{��t�̙���Q>�9s^��k��Zq�a�[��?C�Z?�8u7n]$Vn��Sc�s���1��?��Y��
��hT�"֛����n�'ȱ�x�|OMc��O��FG���`�pt��Nz����Eڈv]�/��IIE7��m6����K���uT<��N*y�Q�rj���:� �(�{Z&��ϻ��8�6M$x�c�w:�g�w��TCJP�Ǯ�Yl���~X���;+p�Vmm	"~_=�c�X��=0�ń�	�c����T��I\����KS�jJz)��ӢސT��52���
�>��Ϣ=F�`u�f��dh�r!� IoZ�X��Mf�Ƒ}��I=�I����-\��X��|�(f��=1"9+0�`��¢�[�}��+g8W6O�ŎG����n�x��t��N�S(48��	&��a��F2�	�(��Io'���բ���Sx�&���D�B2uBё��;ヸ�Z��8UZi�#���;4:�h+��ʮb�;ό.�:1���Lf�Bc�'ˠ�P��a=�r�J$.s�hO�j���鹘��$����=(4�}�M��w&�4�Ot����������x�Re�Ц�+wڻ����,M#B��m׸7�o���/��r�c����E0'�M��sh%%��tMa�t�mݸ;�e����5�
|H�w�[�?��,�������S� C�k$c��*i9���-���c߻������̇�Q֋;U���-�dF��W�&�iw$�eRMt�ڭ,iW�lk�#b��qM�I�mU`��|ުK�����J��2��1��zV�|�!�dCY��B�0��0Letf�`��G,Ѣ��'}�.:��T�좿k���v��N@��#��m#8j������E/�Tg�@g�{w�BWW��?T&v���SX4��.� Vu�qxuj���+AI�ր*�7���/PH�������LL���i�V�a����g�4�� ��~ܑ��@j�+eT���]S��cK�+(0'b,V20��Wiۧ�2_��,|�/�㚦�V��1ޔ���;b�	�rr�:��u>�Y��ct^�36oƲ4 �y�n,
������&bZ���l�Q����3�6o����u�;��������%�0{���2t��F�Ы���'�Զ>P�>x�!��%QnBr�g3���k�reg*���*p4 ��ͅ�m��Ԩ#�a}$�x����΁v����kM���_�w��P�?ߪ 77n���rQ�Nگ���醋�4�����DPTk6��qI:t����_|mTD� �+"ط��ɽ*\�M�,��z�Y�5��:�1�/Z�M=�,�����>��y���bJ]H �Y�6Sx!�J���AU�Bܚ�O[1�t��-����m)1���p�i`nM�,�w�5�W����6��=A�
oSu%��S��xǆ�2N��Q��Џ���%G