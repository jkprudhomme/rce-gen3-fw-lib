XlxV61EB     400     130D9ɛ���l�k����ͦSx�%�܄A���Gνu�Ƈ���U��8��{�מ��^Ls�&�| ����������|CJL����O ����E��Z:��; ��H�9�8��>cR���d�$(0Xe�9S� ���
Fq5��kx2rx�oS��Ѯ�XCm��A��T��0PRSuÅ�7�T(a�3 *�wʬ�j#��/������	��e��wUBm�jv��A�DŴ�;Ġ�o��;�G����`I�S����e�X�CW8�o��vp\,�L>ʭ��mb�%�C-"�����XlxV61EB     400     1d0�>�l��h��[�QH"�y+�*:@���^� ��vS ��OGG�==�Z@���ߏ0op�=��Io)��9��� ,�E���-9:�̌/F���MaDL8����5/�zp>Q�$����l�I�Eש"Th4���Tj���s�Z�J�0�by�B�����H��Ă��:�������1����-0��k�+)R�W��+k�Wٌ��y]q��x�7"&���1\�v˳���,��S�G�2=Ƹ�q��2!�K����6���))]*m���%"�!�XW�j���I�gtt�X�	Ē�k�gi5.���$!6���x
����1��E}�X�
}�c5���R��Ղ$PM��,H;>�I�c��I"\��}�}a���3�EOc3�;_eF���֙��ޜ
�!t�$K����|�M�a��C56��LĮ�� ]�PU��8��c{xp�0W݆WBW���]�i�dXlxV61EB     254     120�vg�Up���GxSv���o��/RVϯ�a���������J�n��~��w;��ݗ�JJ#�
~�llD �w��k�*�U�Abg-{��/}2ͤ�D6�����R��*y����,3��F1Q�Y�yz����W�Tk���1���G�l���rĠi���ߔRfK5��ol��%��Q��;��nK77}y�����F\Ȇ�PX�l\W���_�.p�?*䋙Lc�[�ۑF����DtvN.�֭�}Q���د>�I���P|7��@J�49o�t^�j�E��