XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190���j����#&�+ǘ��U��Xh4��1��;�.A4�P���}��R�H���2�v�I&t�K>���l��d�F�1���`� �霅� Խ��ˎ�5��M-���y>�b��wQ="�*�EU�Y� w������� K$i��<D�a�˂ �2n�oz�p7����$L�N���u��,zU�%TPϊ섾0�kF�Ɏ�]Χa*@����s�NOMKXgy�r�A����):�
�}�2<��%�,�Ԣ�m�6Vt��T��яUW~�tfFPi4�h�������f3Y;ſBe��s��լ�?dW	�(Qt�^�`�l;R��!8]�M_[tfa��|fNJ:}�+���>d���Q�������^i8!��Q�nV͋��ќ=sR%����t�<���4���XlxV61EB     400     170�A��3ڴud����.M���R��Jm������{�Y<ދZ/�ﶅ��5�y|kP	����ݾ&�n�����p
A�T7�R�9?E #�6����#�F�W��݂��WV��BU�S/Z�Z�U�]���o��<fZ�Ѣ>��d��,��瓽�r�s��p5�l�h˨ϼ�eK�_�e;��W}f�9���qHE:�섇���Wl'Y˺�t��W6|��ѸW��o�̭� �L��{J8��P��y� 3$Exu��|�9�$=��뼮��������}O�U!Ǻ�2# Hy��f��vP1�Q+������|�9����������ݚ���1� p{A{�Ȏ�V-`�wlXlxV61EB     400     150�H&�BK�"R0���|����S�M�5�n륕�R6^b�q�Zf6.�H/ J�+�2�8M���҇g�����C�g�Qg�NiB*)�I�Ok��P�Q��rC\���![��Y�q~a�k�ްc�� :U��8@]e�uԘS�-�J-�S#B?an�݀Ng��"΁[���z���z�YgP�ťI]@E��Iv��|�5��?f
�^��Q���#�b��t�[����#)$���F�� �
��~�����H���xT�o�>���.ϊ�R�t�{,���&\!X��� � $��ٗvB��/l_�9�4�����ŏ�Ž���+��. $��nܫM�: $��!IXlxV61EB     400     120A\��*=��s���Qr8{�9��Q�����-��������\���>�0Yh��'9�e�#��N��A���~#@GFh�WX�,��W��:�j^���	@�LN��`�s�\�A;c/_98�(|Xヮ�M9���<7�I�X�%�Ԕ?Ў��6��M��8lvv����3gC򯬵�!d��eL��N����:O��(;�;<�K�1Tg����e�W���{p��`=�'=/����?�&EF��;�m��3Z�9)Uj�<�׺jۺ���DX�3�`@UXlxV61EB     400     130�Ul	P����QOt��+gX����i�rڑT�M0������C��l��|^Yq�R �_�񻌦N��P�����,Ӌ7mʙ�ri$�K�10s�xɣG�S�����d��������\�A�����Q!8�����m��g��?mધ���`���.�<G��9Z��˨�P\z@2��YH~z�rF8�F�Rvc�+|)kP�Ǭ����L������`�o1���s�kPj5��)�G�
�4[�)i�qv&f��^E��_�fItt�(���H���gw_|�B\��K6U-؄t�5�ـޗ��XlxV61EB     400      f0M���F�do�|+p��*���FD�6Z�\=��k`N�i���UQ��.�t:�-ުF�Ķ���3�Ӌ���7����d�r~��=:I&�����O^�'�ob�6r�m6��&�S��?��N��9\��Q��5���6��������WҴwO�I���w��$��������!R�F<�9{����E���
��Qj<
�N�Y�n1pK��ۢIP�/F-����b�|6��C/E�O ��XlxV61EB     400     110�!�tb�5�yC3Oψ6n�pU��]��f �i��q��O��)�C�ϖ'm�1᳐�@�)��\'J���s��h�y�FIn�����'=�l��(���>�k�X�r<�o��ְLD	���QK:$i�����6��)� 韹�O��h�<4�G?�~+��s��=�i*�愑hӞF��G�Dwq�3eg]���b?2�!7M�F�|��A�]p�:����\x�B�ụ�]��o�θ����`w�"�A��H��yC��!scv�E��\ܲ��r�XlxV61EB     400     170��=����J���������sx��&����a'��]0�Ԛ��\�/����N��P��P�D��1�/3(C�-�����An����*g��T��x�/ڋ��赼$m�G�nb�=�J��f�R����������Du�0N�y�9�5��B\�T���6viD4�h)���������l�9��M�Ee"�ױ�<��8+40��xs��!��F�/��3||]Qj����L9V��:�o�~@]��3��1�RRh��s�,�
@�k#�
�7�4� @�9v��A�%�h����-bF����l�4�>�6駯����:�A�8a92+M؏�|r�e֕��||(wBW��]^����W���	pF`XlxV61EB     400     170�G`,��~BF��Zգ��N�?�)��l!Б9,�'2@I]�?��3���N�Ϡ�g���A���d:���T�t2�����R��u�Q��Ej�2ߑ̶$��8U2��F�~�{+�ӂX�O?�܍,����H\��\�¿�h�s�z�]�ǴEuq��}�ϻ̽ P"@�gU��j��IU�v�:F�ʤm���Z�M'iړ`��@�er� ��~0G
��:�}ܩ<�F�y�"}�(1|k4�1��p�$����T��Y/{.��ˡ%��/���Z��Ѱ��{z3ms�]�
�>��3@Z@�6�9e:�tg���F�a��Q�u�ԗ�S��~rg�(�fz�#�%XlxV61EB     36f     1b0��q��ї��	NX�9M�&>0�hA��N���1~��u����4�~+2��'�5��9S��,r��gx#��z�����7��d���?��7�"�8o��R��
F_�-�4?7F@��_Y���%���.r�1��<�
o��\�=�p��[A:��V��Z��ԀkQ��/˫�s��ku1�!�m�(�Xl����N�m�Tr��H��$�/b+�>?\�%�w4��>8e�ߗ2X��AS�ު�(׌��RN�������'=��Bc;�*�C�p yfܔ(LeTy<ܨv���j�y�c'���'ZA]-t����bDy��OT$$��BE#E��Y��nb�����Z��e_ٓ��`l~\y��`˄��C�J�����_��UӖ�Ӹ�M�q�L��5����-����W�������}x'pz���\