XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1804`��٧�/����u�מ�G�/�� �h����e�z��|�=3�w��^��u����2�e��S�k��J�R�������Ǒ%r?����w�m�UT�i��|"�a�����'�W8�\k����DuR`�iFck6�e9��S������S$���UF���+���`��Y�(�?��$����
�D���t��%  [ܟ%��J�[�����_�=�M��w{r���H��
&{�˻c��l�h��2q5�^��kL-:�}*��3 ��B��\��t�9!�f�bx#{x+3�O�1m��&p�OaV�,�]��!|}   ���D��X)6m1�
���A����
�+�Ͷdǈ$U�<��j]�ƙFؒܞ���dXlxV61EB     400      f0=_Ύ!(��lA`�dh��� 	E�xx�؇��C�#"t��ٵz�X;��;��/�A��D�/"�s�i�a�o�Q#��^)g����q�*�}4��Z �7J��i)7�j���2 ����?\�Y���euӭ��T�����6@����V��Ӹ��n��=~���/����nt�۹�yb�i�.I&cˤ5���̯�uG�������0΂(�!�F�^-{Z໦�&�L��Q�#.�KeXlxV61EB     400     1b0�	b+�T��#a�B��	�3�D���O��É��m�V	��+��-&���gƻb�U#��q��e�ܟ6��([�L���2��a�<�d�!>ȮW��F�4(t���[�=Ce���L-���`U
L��F���쾥Y&�>1������	 w����p�Lt0�+��Ud,R�!0,樹8�X R��.�H��,��2��gJlEMB��'�g?XA��lR���=��@��/���!/�ѐ�Nw.�])_3RKA����.`��>`>��/�`��;�d�ҽ���������s�M������^�������i�)9I��֞��u^��%k��q�޷� �.�tU��@�h3V��(r���2��j�<�&{����\T/�g��1{��E��ܼi�E���{]�G*��!��6�Lc�(�'�>XlxV61EB     400     1604[��S�42~k�0��ٛ�.�^�m��N+Q�Z�M��DS.޸F���*�oIut�?Vխ�	��՜z�'?K�d���j�p���Y �^����x'�>�Ϋ.Y�KE/��H�6"H���و�x�Gk18�/MY9�h�L50�ڥ�JS#h�_�U{a�b��Zg�L���q�I��B���nn���.�X���fQ10��B���1��tU=����Z۱���o�l~�v~ۙaGj����=��7k�C�d��3�.��l[����a��gޯ_8yT���M�� 3%L��!Ge�n�Qy�v\������yGW�nV�5��sn)v������6�>��ؙM
�O_��u�XlxV61EB     400     110VU��y	���������"{V���!D�tD�\�?��j�Ɉ��/��������TΊ	�;4���ÖZ�`��2y�^�f��������[�%��^I�ҕ�ւ��B���}��N�L{�F\Al�)6�ݡ�����E9ph(kSA��F�z�:�h���s	�ML�Os��H�ˤ�s�����������!���)������p< ���S/BUH�5��ȇ�?:��*5Ѱ7o��ҋ
	A,��V��B@�3�y#�9%J�,?XlxV61EB     400     1b0*m�yR���+MM����"I�D�&܆��^K�I�l��_!X����~[!XTI�B'�&L�	�^-O��j�g���7�R긧Ǐ�+NI��0��V�N�
�!xpM=�B�:��/e���O�x�"BKv�=�-b�|U��c�7F@>i�+̉�;��G��^����Ȉ�a�����-t�q� �m4ׯ*|�Ę�� ��Z�rF���:(������T��5~�c�+��vՏ]妓Pd�����i{�k$����<��G1
�D��~��vj���sq�S�(]v��ufl�j�P9k̉��;p���H��[l��}���݃ڷ�`��]��/���~���^�
�����`�j��]�J��~�F�I|�	Xl��H7�8����	|&J1I����ű\����fҚ�n�3F;W�]��Z��gC��a6XlxV61EB     400     140[��m<D�E�ƙ�d�؈��,����H*�E����f�� �H�>+�hi�ʻsv��ɈO<٣������*,ޕ�oQ���K�[��W�f��aʨӪ�����div�v�t���M{q�0R���J?/�՟Cc�-����S��-v�W�<�oGn���� h�%��y.�4�V�x�����q9>/TEG��E��<�º�1J�MSM_mV7+v$�A0ce�OmA�j+un��|�y�Z��N�1�����3dDa��!��Cv���F�w�Mߐp���3��	#0��ی���a����S��,�pVp��Ζ�XlxV61EB     400     160��3�r��f�S��]��ƣ,\`n�'�O���D�,��Ė���X9�.QjjF�}�n��'�����3�ѻ_ᄶ��]k����oPH�hk�UZ@��&{�a�g��	�X�����5�mz{7d����ɻ�Q��봢�B��L�&����r����B��eN�*�H6F�z&Kfi�6����APt�m��!
װrG�穰�`pt0_��]���Q�i��vC:�oT��JC��o���S��=5�h��$z��oΒ�|9>�k��5���O@�[>��V#�|g�UG���p{.Y���N���%�W	~�����.R!=|�Ռ��i5�G��d���<�#�K��XlxV61EB     400     190��0Jo[~��*LGKZ�[�<sxÓ�j��]����Z�~��n�N|
�28j�-:-r���2���nT_��p��ҏ�m�H�(��ռMy�MB����M͛㠃��/C9�����Q��ɴ��Lm�І}V�+�|��Z�v�a��n�6R��f}f�������e{4Tc��_q�����J�/�án�1^�f��(c���i�;^�q1���;C5+TW=��_j(0�H=�po�	�D[؉|��MD��ހ���o�C#�]����k�ب�����T�����|f4� ���*������:��I_��TC�ĥy���^[���d�켭�n�N�9�I���m[����*�f�.,R���}'�`9u�`T_1ǦPiQq�}��h�>h��}N#�|�����w�oXlxV61EB     400     190N.+q�vq� ��!�!� ����m�Lj�$��2��h��_�n�F.�VtWɝ�Hd��I��|��ʁ�~�AAM��[H�p����Jt�vS��/�w,>W:f�{���� �]�E���f�DE��Q�S�Va��6�!�4���&����N���t�PeDuw�ǯ�D�����!��uR��8�@1<���4$�s�Z���j?Ғ�$��s�0_n����L�hE�����A��o���≑V�U�qa�Wx���fi�yjb���:[�@h�Ƌy��g��{��� XG���_Aw�W	�ý_��M^fI��Q�I���49������<�@��j���%E-F�d}׫<;2�dC��.z M���2Xp� ty���(|��{��٤���XlxV61EB     400     1c0q*���m`�}�j�4TU|5�h�ܠ���]����zf��7V �~]?r�����n �X^�ǽYA�.p������w�}�ч����L Ko��4�u+C�f������So� ��Cif#�w��s��j�q�\��=Мzq���'߯Y� �����A�"�_��q�,�8����g�59���+1�-�/�;��
eB27��� �'�0j��<R�9��An��7����i�E{�Dp����������tW�QO�yat�_%����j3a!���GCp�шE3h�J*�.;	T��5����e~M�9p@nm��� A�����s��Weڃs\Z�#G��E�\�7�m�O��������[!���Ջ��c�94_��z�1�o�xԲE���׎��� *�1>d���LJ���ʎ������8�[��9zXlxV61EB     281     100�Ǎ�:g��;��jm�p�0��C��`��M��5���1S��U��,�/�n��o7܃/�����e:4�POsz
�0*�c͑�����Ny�n �"�Iv��;܊�d�K��=��T�Q��xbyL��X��7p���T�y��|����F�k�R'�hz��aEx�apf��jx!C�2�I��7�c���ܯm�:��q��Du��@�cAC��������j�s+7�}xE?�F~��8��\��=$�v��2�r ���k��-