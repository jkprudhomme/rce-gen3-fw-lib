XlxV64EB    15da     890��=���0�i#^�:o�x�ˬ�Y廗������r�1�*j�6K������O<"�-)׹'AqQ�pC*̀cz�Æ9l� �]xK Ȳ����|�Ms(g��r9��ӈ04��-,[d�/����p%gk,4��Z��y&�W�"Tj�`
��s��?)��=��~��B#���{	>��$_�,Ӌ�m����<ф&�A��ǧb��7n�C�>�T��l""��I6�E<`������+���\��&�q��%2퉘v�&��3|���]e�:e���I��yĬf�]O�P�2c
g���꽁�e��T�'Jm.18� l*Im�&��	E#�����dϏs�'�/F2��'�i�`�	m8%e="��$y��;����d�JL�������Tt��2�@����zU\^��X�oƼ� ���������c)� �zq�+��7���H�t��Eِ8�6Pb���zd��\�.ޅS�5�Ru��� ��V���Ǟ�G���\i�����O<1����X �V���]Q��	̃��z��jod�:0]͸��B���,/^��9����ԍ���*�Pƞe����#�!�Ctk*3�Bi���j���r�_������u��:����V���	�[�D��fm�dF@�t���F9[�`�@��� R�M�u�6�d�����ds���Ȉ
�]�C����K�®qf��Wj@���"�~�_̸�/�}�P|/pӤ�(�v%����q��L�����/�{~*�� �ۄ�BO���l>�F4 �\Z��ӌ�H�%A�"�B�n/����ƨ�7z�t`�:�o��-E1�~���z�A�J�L ����-�)1�ӟB�Q��qR{[l�B�V��u��Ex����+.�л`6�=��,�\/D���4����Dx� s1��ZPֆq�97�<a�|�A��S݇))4��d)Fh�GG2nq��&��:��C8�M�о*�v*
�cJ�u|T�O�
͐�{���#�d�O�B#ބV6�xܳ6��"^�[b��1L|�A$?>�rw@��t\�QjZ�yQO�l�\�?��[8��CpϤJ� ���"��3[,x<<q�5��4�D�i�8��m���=���D�{w�TUqOjS{ጊ�r��Y��(.0;����.�2@|�������,$v�������P:,�^������ߵ�%g�$����]��A"I���Z,�)���uut@qa�~�3R�(�?���C�̐nk?�M��`j�ϯ7c3�,E|��V�/� �l�T+���
�	������]N�<��{��9��$����Ie�3�'�'�Oᔸj�u\�h��Mķ���/&o�(H`�o]P`��'��d~�)<l�@��������IS}3���#������Oс�M3�Y1u�H�O�h�/�S:C��]�[�i?�@b�06��&�!�k��^�Z8�	L��5ٍn��9g��B���p��^�T%�f�^4.�/���I���9����	���݃v���	�=�HF:�Ȇ=Z%*4��k/^CX�e��T+U7=%:�q$jT���Z�C�ǝ�]�lO]���-�PY��f�_��Ũ�'豯�����1x"6�]�+o@3�JE`�'�\�BO9+��emDY���~����"W�v��ۛVcM�i����.�������2��F�
=��x�����k��	�iN9����#�8P�#�wr7[?�������/̋1X�Ύ�O�����xxZ#�~�1>�Ʀ���y��x�����LT��۞��B��7��S
�?���a�Zÿ��aF��!�xR�&�Q�?	��
�SB�p4
3��#�d��/@�ޢ9���+�c�/�<Q��{�zy��p?�_�����^����ʪn��5/؈�P�r%ȄPF��d�{6�	Ҩ�o$���XD�5��c93�'�3���OΨW��OJZ+����M�S���n6�X]���+�h5��y���^��~փ@�O���x޴$��K��ٙ����<T�P�rs9T�!SZkq�l8&�?]��c2˷�ST��̪�02��4v�u���U
���5YJ"CGv�X���b_�حR^YUDz3;��X�'�Sg��a)�m���dT8��FĐ	�p�