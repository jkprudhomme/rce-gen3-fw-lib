XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     140d�9��o q��-�MR��7$�>`�%������.Jl�!,V)��M>eFg��A^���/
�GNx���p�c0y����ml�Q�%�&�=�wK���E43��L�?'�f�F]���*��.���<z=;����~��~�дJf�@�5T�Bn�}p�3$��mh��]���ٸ��$q\�� �)��=Y�ԗ!�B�Y����%֤�ݟ��Ⱥw���N���aW�
K|�i.��ۓ��v	�~�|@ZHK�M"9>���m{�P�d�'�c�6p!0��1zPt����U�q*��W�U���B1����XlxV61EB     400     160̶����	q���C��ʓċW)�.9�j)�֯��AL�,<�S�H��×N���0�,�5���|B�?��;��'����
��jyNr.�	,�"�9R`�[����9�'7�Z����&2g���y��y���4p#���M�B�h��S��:�'�<V
r���� Pjd�Ԁ��~��2VHV�G��Q���U�6�_
��#�=Ĺ��ق���4�QTa$�s���W�8��c4�ٝ���JUD�-�:��l���%���3��4�7�ۜ3�o�����D\y�
��=A��_#j�U���2I��-]�cJ.Rf_�S�~��1`��O��r����E
���Oem�D�XlxV61EB     400      e0�&���t"��Y�7����<%��uf���dQ֩_r�Z�����nٺք�۬�ȹ\�,_�y�_�r:J�:e<�Xp��[�/ �w/v�o��e���U.��o�V����❈�[L��o�x����c���⫌��c� �m��\�r�?��O�뾝���6`���LQ=�s�1�&u�դ�@�Q��ݷ��V
6zך��Q���A��<�����|��XlxV61EB     400     120~.��� L{�9��DP�����L�[�l��v���f��G�烋���4��� "��e#3�t�WyJK��w,7T�:�OG� @�S�Ubbs�����cJ�
8ǎu`�\L�`�|��-'���L]����ZI_���u3^F�p��cX�%��N�����^����O%��|��)Ƅ[�(8.�b��M"�*O�>�Y����w��T�E(g��-����Ω�?���n�_�kz�p��9������5E�?�g�yE"��ȥ	�'XlxV61EB     400     160���y�.[�������\�$�ɽ7�̾�'�N�:���n��G�7,�I���g��+�d�N3�S��B��d�t�a'�>5�貿_�k`���H�l&0t�/TZ%��`Mf?��=o,�xf���̛=�Vے
@n��0���c"�q��o(�R'�+�!c�������2�
%�1�1Vf��&��UG%�Qr��Q�5(�q�y�@�4�g�U�X+�2�_% �����|U�C� ���flB�¢|�A�3�Ϝ��^��)��S�ӑ�/��(�g�$�SR��^
���ږ�%�0�����qMʺ�x���m��hcg��q8W_Aq�{$XlxV61EB     400     150W����c�eF&��ţ�M�ma���g�\C@�=�W�@Y��e�Z%"N�o�Q�!���x���c�t�N��qi�ԧ餳Yi��j҇�g�� �q�|���{jy����ZmY"������ }֦d~��3R}� �L�����������%/~B�]��FQ�x�=��7�?LKۊ�֧���2�|��Ik*WI��[�]x�Ϻ(Rj1Fōl|���*���ף�
��<��G�\��x0��@Lك]�%T�YV.��>��/P�"�Ì#m �/�|
xg�kx�̼SO�f�-;�&�`e�G�U�1V��,2�:��"�ɥt�q0XlxV61EB     400      f0F�)=�� �}��iP��$��NV��*�'���i�ķ&�b���7$��C���`Whߍ�F��E�R7���
�>Z�̄i ��i@���}+Yd�k\@_f�h�	��,�~榩�a�Z�JK���Lt^^*�-�i_��$��4ރ/�p��7,���S�0`ϻM �mY0�{e�&sX��;%[����Y��o�u��i���V�*�g�`�3_��y�th��nXlxV61EB     400     160�vݙn�}�I�#0M�׀�]A�ƃ'����I����F�镜"	Y[4G'��}%=ϩP�� ]���xd��Pc�+Y	~�wB&�y�'cҦ�>g�]���a��|���M�����h��.�k}F��,��*"�,����{�X�Ѣc$ЄU�(gǩǧ�������{csf܁c�W�
�n朹SY�[[ �$I~c��`������E���7�e�E&�`zK���H*&�!x��%�
��!��8����ҿۇ4o�^�f�Us)�`�D��3���D#s�=Y�D�qT�-D^����AL�N��S�߆Z.-�����<OU�@Xxm�"�l�������XlxV61EB     400     180͜�Vy�ovn,ۃ��k��q��9��ľ� dڡ;� �ŭ�����lAZ�Gc��۸�IxV�3Pf��F�n����P9m��R��S� �S����+l�ƴ��̻Ϊz��&�P :UłA2H؍���O�b�c9qoarG"�A������j|Y����0|������t�U�C��N��L��ϴ)l?./��)�*+�'3��^��WT��;�5k����������(����'V�N���������.Rn��;z�NC������7y-�_���+m������m�I;��/�`���/?��{dI��)i�؆�t�Ŭ����}�� �*bB4pSN/��Q���>G<V\���N�A5l����FE� n�;�Å�z�
��O�K�XlxV61EB     400     100��4o��A��Y,`;fܘ�◇F*-�ck��>�*S�S)����R�7_;���oW�xj��Z
�tg�`�9�v�Ok4�1^����{y�Բ����!	���Iz�3V�T�R�-3!��-�mb�J���*���=<M�7�ѩT"?����C�o<�����qq��|�s�a9�=��9r���Z�0�}�K�.5k<-X���}�?�{���P�sٚ3aFP�8ل5ﵔ�?{R������C-�li]?�<�XlxV61EB     400     170(efgc���P�+9}C�0Ot"B�n11/WG���S
��"[��q9��7�I1��t��.W��w:���>j�~i5[�xRe��ɔĆZ;��эW�����q��~����F�z�y����|*q[,W{,c�n7m@D.~ʦ��5��o!���DH,�C��Ʃ�W)}�:�Z?W��ٍ�����c�`�������4�>Ǣ���p説���--�[�aq��8�����Q?���Y�|oe��h۪�]�q^o�Q| Z�j��1C3��0[�^uK��^��c��<��{Q��=�3,yi6c��^��wZ^>����^[�յ��9p��j@<��3
��L��$f�<�����!�*)�/2�|������XlxV61EB     1a6      d0��x��ޢ}W ��v����ۙ!<��� ��
x�����ײ��e=��U}G�Y#��>|�Yʘ����*�;	#�h�.��.O���l3�/�塄�J����k-�U�Ȫ�9mfi��ݷN"����6���ǀ��C=t�� ����,���q"��J�c3/����Uob=�O�\{]@�H�C��,uS��	���8ڑk�e