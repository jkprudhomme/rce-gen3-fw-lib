XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170�@�b�����-ؠ� 
!#?��X��T�X��m�-d��� س�FM̚ä~�o�q���N���T	�p��`�5z����W�}�݊��l�ҷ=ƼӦ��Ԁ.�k�rL_�|3��v�#���Z������_��WQ@�hP.p��|�g� I�<�{	c�4�1�Q���N��ըd�Z�$#�	dvI����C�{Bw����{��Kk�K�)C���Ȇv�>��K\r��,�6��T��Hd�*JM��i����T5EcxW~LX:����Uŀ���]��-�]�.�p�[����I�wL#@^���l4�#;��"p4<�br�H�%O@��,�����QttM���U��'G��Rc%1XlxV61EB     400     1a0A%��2�D�Z�+K>�����tɫN�YJ�9�6���G�t����8sL,����o��>�3�����.��a����O���8�4�m�
�7_-;�Γ\��?�Zʕ��0�P�p���o]<����\7q�!�w��^H-��o	�h\��p�8�_?
fl%����dk���ˊ���X�kt��
�	C�l g랥`G�$a��	��4��$t*@V���kl�з��@��1Z\ޞ^���$�*~�yu���E������+ᒼ3P%񇫂�qʂo@��#��C���4~B*�s�F�y�f���1Y,W�}	�V�j�6�]��θ�����pg�� )S�]��{�Qjh�(/a�j���:�1Br�t$N3�T�~�eH�x��K�H���C��Q��O��U��3�XlxV61EB     400     1405x��Y�t łh�۹�mV�H�+�m�r�A���! ��&!R��C9��vj��T-�ǡt�&�p�;���9YC˷��~!yJ�#
!l��7�E#&�^�	���j(�=3� �k�5S���)�ael6T�5�k;�Z�$��41C�e�2yL;��3#�����	c��Y�uU0�
�t����Z�m���s4�t��k����o��*�v�i�KR��T��ߥ�n�+j�:��ʧB���-Vx"��0(O�/U��BK.2��q/�*��)�4�����x��#�����ib���x�|�]g�ʠ:en���m#dm�XlxV61EB     400     150�Y5��FJ��?[ֆ-kh{�n�}q�Ҩk�:��0�	S�_/�F@j��XD,���۾�(�Wפ���N��	vYJkf��]�1C�c����W�㼎E�l�d`Ό0w��c�{�r�#���;��M�����Ѭ��U:������ZETv↤��&Ȃ��5��F ��Ξ�ZH�mK�6
���l�H�ų��Q�XQ( mstF7>�l:��/D9������ƠHK�g�eSq���<�U���5��O����@$���!�f����;����3���C����k��cqi|yk{��LL��������e�q\�@�Q���rA�+XlxV61EB     400     150�j,SF!��nZM�b;-��S�f�L��ۗ%@�K,�;AG�p�&/]��5�Ѽ�~��(J]�5���'-�x�6Ӏ�
zƶ��u��T5vseQW�M��^͇¼���3����q�J��(I��;�J %��)��2@Q)�q/ld�!~�W�Y�5�Ӛf�}��u;	�C��钓�~o�:o
�E#$ ��6��v�Yl�d�ތ�3��m�a��+!t�ȣ�??��+�:aY�u�A�S��l��n�3��ev{��#PBZ@��a���Kn�lr���AwBm�]j�z/��l�6K��g���5"�HF��Wy��)8��:-R�u������d*XlxV61EB     400     150&#k�!���Զ�(?�ۚ���o"@���@��{j֔:�W�f0�g}..�T��j��}�:Z\a:4'����u\��6��)�@2=�{F��Hxv��:�n�E�l��Pg����5�P��|��HU�|��-.r������)�2��q��,7h��>��ˁ؎[0�K��Ԗ6ϻ�R�DZe=g�x�3޻�'Iv��_�����HfOu)��,��xwM�,�#�X��ay�_[x�����a()ڵF�nF���p%\)�d4�<�{�W',�"�2�2��-Ki�{�ׂ���IZ�80�G,��Kg�[�UEq�{�3�i�ߪ�R�[2XlxV61EB     179      c0��Q�n%b�]�튼��6�E*��]������H�7aPU�n��×T���z�io�*���~�]
��Y��ުp2=�7�d���SG�"�������Ξ�u�Ũ��21'�+�Y��	o̅X�ttN)��f�&��oy��S5��+�.������Tu���e�^Ǌ�4����O�S��Ҕ�H$�