XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     190j���ړ���:����Ծ8O
�lM�_D5vb6&4]�uTY�-�����C�N��Y�N���2�Jk��+�%r ����+go��j���T��P���y6Y�2��Fd)U,�CՏ��ZoH��9;�+�~�6h{��:�����S�'�>(S�]C�H@���P����+64X7�#���#��0��V�x}���O�P��/�gӪ������O�yj�d[W]�o��!���x�=ޱ��]M�q�t�}m� ���G�s/�U�|U����3�J<�cs��D�C(�̐nW#q��_.T��W�,��vn���8�u�9$߁��e���?m��|���&�O�knK��S�z$˫�~Rj�tb������F�m�Y���z�+C���mL�񚀬����N��00 ����XlxV61EB     400     150"][���~1(��tB6��nZ�%���n��q�bӮ5|�rH!�Q���2a>2��HB�j��)0�!A��j��� �^�a�<֡��\1�����d`�9���y���ɺ��,G�8����H���۩����¦;┯�s=��$\p(;����%A� ���e�lBJ�d�)���8�@��(z���4�d�Ea	x5�􃌀������j�m?a���~��p�0�\��:��t4�I�(�:(4r	^M3_TpS��z��v�E�l���!�'�s-Q�\_����TDJ-����oO�>B7��r���>_1��q�y.dH2��9�1�t�l�&���D�XlxV61EB     400     160�2���>��lQ�Þ�(��*R���u��
�-uo蠍<�&�\9������U�-���n��Jv�n� [���.�^�����!a�QW�C�$�CP��<��à��Iv�Yj��n)�	b⅐��h;$�A,�ķy���<�>A�\f�آ��/շs�˜���r���\	2�'L��Z�g�Ғ�T	���b�-w������ͦr>c��H3HN,��E�bE�=���(ʻ�K8;"Tr�g[�\�����D���$5����
�9�����`�K\��A�#�]:�����
W���Akx;6��`-������Ƶ�R;UWG�c��wl���V$yQ��WXlxV61EB     400      b0�"L�����%�!]�/�8�	`m��2�A�D����1ja�j����x��,݁��3bmVɼ�N����"�@�#ۃ�BUs}�T�ڬ���N	����	7x��牘j��G�?������1�;�:L�,x�̚7)���/���?q�2��f|�Ϭ�!̼��(�ws��鰍�������,XlxV61EB     400     130��C�0���iC��goM�SG0��O�����|���r|��N��_c��#��_��hRExܩ`��n��yK\D�G��b���P�3�ʪ�n(BQ�<ݑD1l�\v�W�c����|�V��w�ne�xT�G]�|�]D�3s��o���v[%I�T��b[�ƭk��gU�lxW����H���ܬ��$�����ÉO�A̐�3�R�Ѧ闍c��*�!8xIi�kC��o��mR?���|���La������9B)c}�B^-5%�D��~��M'~l~ ����+�]f�,���nXlxV61EB     400      e0o��=�嗸���	�:w�E���xhF�$��c����҃�_)����V��ˆ�6J�ۖ?:<�7������e�C�����r�u΂�W��:�F-��r��[��M�ki�A�0'�Vz[��Zj$;t$�!�Ο��}5���|>(�٩%J4wE���A�,߸no
�mν���(�{K��?���?O�<A}
�c�/P��y��Yi�m�XlxV61EB     400      b0�x��9eʵ�Q��(q����Pb�f�P�mʗ��v9ɮ6�U�smG4��Tc����w �b�pn��{1�(%`P��<��P&')`]����,h?,�Y_VgN�}p�7| _�~�0)��y���Y�X+hIp�3�"� �2�T/����O��X�3��v�B֓���K�XlxV61EB     400     160�]�����L��x����nEQkg]kfus�����)��Q_8�+�_t=+�����K��P�l���}�Y� Х!�&l���?BȄ�9�q��9͓���8�;/�����A����Qy�wRC/<�Z�+�y��I��f�mzW���}��D�+�臇}�����@Q4NQ_1���lX4S��5�ɒ )�����c���������my��|2�>�4�7��]�w�YT��JO�(�g�"M�9��	�g�p�;;=q�'`"���pU���{&Q���e��D}lt�(��QmgH�>����j�5���A�1���V|x�ц/W��n�����3�������b�7�sf��XlxV61EB     400      b0�,ɡ!�&sΛpfA�8+}�r1�Z���o]�=���U���(f�r��d�~���}�R
�=4	��2bw�o�h�� @�Zq�h��B�,��S�����_�U��sb��?��tf��⾺M���:�35.`Թ���;�-M�4��O ��:V�脏�(}Ϝ��5��Ի XlxV61EB     400     150�C�?���Y�i�,�A�G�y����$��h"�\W�R�����*���{=<Hu�!G����.�����+ۉ���N]�y�@&�س���i�̡+�2����^�tXSD�s�+0�B��?$z�2��6w���G���.��u�̏#�9�"���`�er�����qЅ2��5T�kZ9������&�n�6Y?��K~� ��r��HsĎƈ(XE-�?�'�xk��&7Y/cz�@U��;�b}�;�YFȽ����Qv.���LJ����i기�r�ϰ�ye3�ׂ��Q[[������n���X��� �py��x`�HR�SB��b�XlxV61EB     400      d0����񓜬҉�1|���ˍ��&��-G�}�N%uc/��(���A�K�2��>���3�� @�Q�F{chO����m�i{�J�A3b�ts1�0�6�JկM]� _jPw|�J�^���:tz:�Dݍ%�����\�+5��J*<D��rj�ª:��_��8>������Md��F$��,.P�Ѩi:B�.Z���3��~���e/��XlxV61EB     400      b0e�6~>D���3[�]�c����������g��X�ly��-l(Ē�!ht��X��4���I_�50�:.<���&�� 5� 2�q��=��TF= .'o�u,��U���\0go&��fe?��!X�M�:�s��b k��رؗ2Y����+
%�z<N2��^��*y�x��}�XlxV61EB     400     1c0�N;���Yf�E�ib�������0�#�b�x��Z�E�wf迲G5�����d����=&��I���~X%�fL�E+�n�����uE���&�Ŗ�z�[�>�X&�
�W+���W�� ����N�NQ����,����u\��<v����l�n�X���S��E��ElS�j�z�� ��r�.}s?�Nh�B�3���R���}<B�Q���޵�3W+
�i���l�р�H�{���$9�Z@���nc=R�Wu�l<l��Ƙ���To6�I5�?����3�4>$���o��^H��	b�0�����cu8�L�%�L�u��b{�[vV@pX� ���-/mS�Q���[ˉ�ʋ_��uq8%��<G`r��B�FC�(J�/98q�䐵��w�����|�J��bAPD@ap��(�~/Go	%ֿ��d�y�gN�,o�'s�!��?�XlxV61EB     400     150�s��t��@�ʭ������Б�(���e�:Puy��7	0������zҋ2�@P�E�d��iq�٥�n�uU/!!�l)���{�i��6��Yp8\L�b�"���¼�d�����6;4sM�UDF��՟N�����G�j��("s�ʯ�]8[I�P�g�G���# �?P#Z�"ݐw����%q�5L�E|=s���`A{+�xQ����\(B&M�����|���?�n��.��T�VڳG -��N���oF�t��T�3c�*��[������i�Wu~����=�~�,m��P���+a��Nh�"����c�J$�fS5�]|i| �f��7\�*��XlxV61EB     400      b0�x��9eʵ�Q��(q��1��b-RYǌ: 3+-��*u���q�T
�|cR�0p�L�4L�$ͬA)6TY�Y9��gbg�ʍk�����?vs��@���%���A�x��\�Rg�7�ѯ[`Ů�d�4&���G\?D4s���:�K� ;f�*��_��F/m�d�
�� \�k��-m5+tXlxV61EB     400     150��"| ܯ�lOGҧ&3����9s�Rp�y��!�[��SŤ����q�5�P�=�y�����f�ju^��G�Xz�c��d5�P��v�@5�\�m(+�kX?1��3n-,e1����+�~T�WΪ�n?��;����E:v�SF��vy�j�D$�97}�ǝZ��9P�B٣{m\�H�Ӹ�E0�K�8=[����y��g����^�il7�+'7fqe�!?.�W���{�]ɺ��>�^����}��An�C/��aewsj�4e��/�e$#�T��Q��V������I@�H����UH��W�j�S=E���o����p����t�w�XlxV61EB     400      b0�P�����υH���X99Ӎmۮob�2��J��O�F@!i�g�/T�7�_��jui���)}x�����f{M.:=���Dj�5G��gzz�x)�(�#D�-���r�"���)������$������$���)0R�7aĂ��h��D���C%��1rJ����JXlxV61EB     400     100���O;FJT�>��?2k�o#w?�0�')	c���|J,{��8$8A��;P���L�a�r^:��m}����q?^Bs^=	�����0���oL���K�'L���8.�H��+�\Z�P<��������!n O/�e�Ѕ����4���#�h���U�w��O����s�x!�zO���z�X�ʆ��T���q+G/ȏ������{p����-�
BGXKq���?��S�;s������&\ŐH�R�Ū8௫W
���XlxV61EB     400     120�T��@U�ɱ��e��v���Q��%¬��~�_��>�Z���k�g���pu�f��ĉD���I�jg�w������8�T��-��}Ͼ$��Hg��?,�Q�6�OƾMT[�$,x��@�' �����5}�&F]��,/@<����(s>~<��������;���a(�����읨L}�	�le��r�������aU���N�]wˊ��k�k�xn�V�s%��|�;n,��>zb:ߛQ#��6�~�`Q�2���V���`ZX�"���x	�0b���RDh�N��XlxV61EB     400      b0�Bs���./��'@t���$"�3j9�bl��v�]���?Ts"�����������qt-����*��)�𲖲ҿ�n�U���t�n�������x����u5h=)��C�,k��`�O舵#M��N�7.ך��T��@!�z�M�R���[*Q�\[�`�`XlxV61EB     400     160ė�<,�w��OϾ�-�����%_�,��+L~K������B#"�(~�|��;d>�Uug##y�����e��D�y�sJ[��ŏ9+\)�iڣD�N|%��,�_�:<��db�+��8���4mQǕ\��PVkfWa)aGx(q�*G.I?�m���hf�u#_F[i��'��G�fZE�����ߢ#����r����c�������C(n[Ǯ��wXE'�M|blf<>b��R��"���"�%�l�*"K�Z�W�&�a�>E�qI���4a�v�I�]���>���w'�����X@&�m��6|�n��q kP�$N!�m4C�d������7�D����XlxV61EB     400      b0���z�� ������A�����ly#�`�X"��o{z�c/���(�~���C)�p�v8��[c����
��LE��/�PX�F?PUIL3eY:B��<���Z���zI~�J>�����RJ�/��@gk�f��c�>z7��-N�~�лib�_m��4����EXlxV61EB     400     130Td;�Ƅ^�݁M16`�Z��2�)",���Q�K��>�%�*"��� >��s"ߊ[gAޕϑ{��M"0�����U�g�L�CH.5�բѶ�9ȿ�:�~��4y�-��t�Yk�ㆍ#�›p���\B�ҫ9~.VWb�4$>A�ms�7]�
~�����C{,�Y/V��a����}�mЈr�U�t��]��:mE$i�'�M�@��߀e���o�
��:��&wֱy�:&�x��rP,�GuI�����	��D$�e�l��M��;EYoG�$�	�7�J@�⫾L��ᓔ%Wi��C[XlxV61EB     400     190�eK+V<��7P�v������W��A<�z��/s�m�	k�[|��v<�#��b򕀮�s%�oܪ�{��	�lc4�UNzw1PXbf�����䷲���< ��t����}*���HfS�/ٵ��`8�գ�ےy&[
9�A�.��Q��8AS���:�4kUp��4�!3��I`EP|������(��+����B��x3��dʼv�Wk�2�t2s
�h�X�>cS��&q5� ���&f��?�w�V+bXL7�	���\M-��c�}�F:yfȂ,��	� �˪�$����k�����L�� ��[�hG;5~��RQ��g�����[[�	�.t�����k=���f�a�q6���E�mA�Q��2��ɉ2�vk��XlxV61EB     400      b0�P�����υ�'���l�� �l�*�^x����!���4��Ű,��RY'��x3��Q�`�4���e�.3���3��PE>�Ӿw v@�I�@eѺDY@�si,���qA���Jb.J�N�hh�H`�H{	�ó8�Bj�ot�S�|�	���rvW^�%�X�XlxV61EB     400     110ճa��������}E��G��
e�J�<�XBd�D��m�������ͺ��_ʉ�yS��I���/c��V+�]��\!j	j�sF�"9�<r
� ��NsA��<��h��@�A�e��|�]�1~�
�s(�pĮ"#��+K,n��L�J�n��P@���PK���^MȂ�T��5 ����X#��<�EF����F�|zo������d ���=����E3��U�i��/bD�)���G�����!��4�/�� ��d�ǉsκ�d�%gXlxV61EB     400     100�I_�G��k8�b��~�a�S�Y�k�������r7��ܪ��!�k2Av�j���ʕ�����`*�A$����=�Y��L�~�S��E����������m���*L�62�Q?���H�K���O���a����sP�)����|D��&�曒i�6��uh<��Z�q��O��nN�(2nj���k�F>mxo��*I���_(������{��٣��:��֚( �?U[��8Ȳ��;�=?���XlxV61EB     400      b0�D�ȣ�^�׵�I�F���q�B�[sVy·e|�`���a1a-�4l�v��;e�P�gn�A���q�x(�2��5o��0)}(ڒ���ݫ3�	�U���O�񳼊WOQ���鈦�Ļ�<G爚�#:1�r�u���IT@ר��YB�m���gv��M���j-�h{�hIr�ݍGXlxV61EB     400     160��4NoV��;�"<��B$�=�x�����o�%ϭ�u��\L�ҋ�: jzkAC�ߴC�������(����`);��HG,K���)�u���c��P1^<h�����q%��n��F�⛸�g�%B�b���j'���:;(:�i
�m�H���KV�s���w�����[�~�@^�/@u��,�}�wΪ��|��P�S��bD�d���0�\ӂ.��]���ݐ�w�V�غ����`�����vI�E�i#ٲDQ��Mk	�/�/6:ų�b�
Ĺd�ʏh�x����k'�������Q?��?���2p�~�T�T��r\���x���3��T��U)XlxV61EB     400      b0�����l�+VR����WP֟XX���M��������$`(��&�-��;�H�i[����?k�[���W���|�ra�07�����BMoo;���M��
���p�6/&;v�	�GTpXI(b�ug%(M}�R��M�@34%�ƚ�K��lj�qP
�8��L�5c?�<�!�XlxV61EB     400     160��ؾ96�#��瘠��&��k2��E�B��VCC��}L��+�=�.�Sqq�O�Kĵ)-6]s�L��U����,�8hG0;P��Ɗ�[��H� �$�:�����R����込��t�t�TP�������?����E̚�)����P�H�ClJl �,F������1�r�u���4�#�������82I�Γ��n*�R�q��Q��b��no��A�vʕ��&4L��Y"zN�g�Z��6��U��q���k��=����ͥX� w,��
���8�����*�����}\|1(�>�C��H7iU��
��K `ίZ�ZZ�ח���
�gտ�}�V�XlxV61EB     400      b0�h��k*�s1�#�w���w1�\ܼ^a-������l<>;�]���L���6`������C���L]�֊�Z}]�|̃�(8��	�k?"�ʃ������{��׷��p�N��kC���^�ږ���3�Jة��� 9�*��1��������0$�@I�&)��L���-C\��dXlxV61EB     400      b03��������<�TM���)Ӑ�7�S#gl�֞A�L���;�Q�ҕ��,���ͬ%���8I�<�W��ܵ�����ŕ�d��� �����$���
�3:5�[E��B�R�Z��	Ѩ�cC�}J��B�o��KCT_(�C+�M�@І��*����>m�K�Vo��XlxV61EB     400     1d0u�{��Z��~�ӿi�Y��Ѽe8�Z�T����%4���0�(�˜;"��h���U��cp=��Fi!/����:PK8/�@��}�n'ws[���C�eB-�C��[b=�%�wlCX��%�b��)|�/�w�խLАE��U~�fQ���|��Ϻ�?�3���xטd)i�,yu3���Tl��$��!4�F���`�)�8������.��^�6i��dG�\6�p��&��L�hpwZ�FO2�����U�Uݟ��e.��g��;�w�^��e>�I�������Fɇ��G���UZ�7�i�
�XY;�Qd΂�b��f´��LE� ����j�G��P�.�f�O,��`�/��m���!�����}*�j�W;͢��!��<����4
5��#�حYq�A��[<cHD����o>(�L�ϲ�j��G���r�@XlxV61EB     400      b0��k"aA�oj��2��ũm�s��=�W	����/�s��v��)��D��)uc����ijX��Q2�z�^���LJfd8�d�F��@`}:�e
�I[����&t��\�Q�i���+h�0�Qdi�BKV�·f�<9��&���� ?�;'y�<X�R�Q�r�&�=A�_���bpXXlxV61EB     400      b0�^m��C]������
���p����M4&~�b��鄑.��ǌU��X+�o�/R�.݅��[vt � G�jV
�Il�6tR���_%4�+�U6��{�8]zS�M0Z'��1���n�A�J�����R$g�{�?ڕI�륋A�]��I��RldH��(��"kR��XlxV61EB     400     150�rG/D�yB5?���DD+V	�"\L�:�u�w� ��>�ԫH�?�<�*г�n6f=20Z��(�gR
�Է�e}��b�G�K��f��Q��N9v�(z�L���#��C���R����h�,��X���4��L�k(���ꬑ�q�m�T �F��8����(2)�uC�3�(�{p��2�א����ɼC���t���9�V�p��=M{�������c�qEh��>�dR��>�K�,?��EOͼ���� �ч�S #	E��v�~4.Ѳ����v$j�qq�Zj_��6A���V���ɧ^���*��wu��=�-0�c��W��R���XlxV61EB     400      b0�҂u��7�Y�Uk���T1
�R7���+�S�v<&����,`?�nl�+��p
'Og����G���/�Lw1����}r8��Hm<�!���Y'�yA�!���50엪/꫱;� Ӥ��(�rl d�<J7��+��� ��� &�4
ƣ<�>@R�L��5�P��I_XlxV61EB     400     1808I)�5g���Q`4RuB��|[\�~�Qꡍ���è0_n1*ЍRH��ԫ.�!�[S��J��ݶЛI'Tu�N��).��]ܳ3|foC-:sYͥ�5tYb�pM�	%��Y[`7IB��L/}��ʆ��j�|j����	x�@��_��o��5g��n�V^�Դԇ�ڻ�K ;��؁��)�D��ss��!�Q�
z_������6��#�M}�S��Ƞrn�Z��q�)}>j����9���B����9�
��B�jc�TV��%@85���84���f�KB�Q�} 6��ofc�$)N� -�+��}����H{�|f�G<���!r7n|���5���I����הs�K�������$��o�XlxV61EB     400     130�Y���z�g���icE�f櫓Lu#hЉ�T:l5��8�����N�*@���sT�g��3��G!tޖ{+��<ĕ������<�i�W���%֙�H:ּ�P
ܞ@������"�ӕ��ut���-p�4%�ך�Ȳ":���ϕ�́�ت�*)Rt��
��1�:|�����{�P��$��?�Y�%&�O㼾Tјoyxr&��K]4%)��	��z\C	BʥO	@ɀk��fB�վ����U3�P��Ͽe{C!�!��y�47	�u�2ʁ�&-�Q^F��	����n�S{-�XlxV61EB     400      b0���(|�U9�<�E�K<�xDQ�\��lCd �
��G��@|z�Fu�v��S�� (b�a���*�Xa]�F���bN){�!���Ba��a�����	n}�������q_.8�*�y���rw�MR8C��}��22�ٶ?��=�3�)�	���q�uĒj,��彻�Y�XlxV61EB     400     150��#4y�;s춓�t$���;x�Q��!D�Z��5'˝;-q��h]dRG�K�z Wl�_��.R�� tgJ�At�����ʗ<�At���Վ�6�3���-d�>��NЛ��������m��a̧d�;?i���-۾-����qj�VD�ȣi�jV�=� dH"σ�6�!�DOİ�l�Ht��p�F㌷��Db���N�b���M��ܺ�=,͏���Cy��ȡ��h{�`��,`uʒgE>(y�GS0l�	X���?��� f֟+Z�=�6J[� :�`&FX�u��E��9��������:dƪh��z����eC4-�J]?B	�54)�LXlxV61EB     400      b0�h��k*�s1�#�w�	X�����!��&F����=k��\���>�/ �	���{�PZy?�=�F!�'�V�!�U�t�I��ukח�l���<�+� ��PH�<��1�3�6c��
v����_��\'�v�`���.)��By�V�䧲ҳ'���/�l/,
O{�7���b�}XlxV61EB     400      b0����%5�^Vd���Se?�Gm���v�1{=���$ͧ�
Aon��s_���pb���V�H1@�I��I$�?pK���ۼ�ێ����햲M��j�a��V ��a��k��B�m�Mǭȏ��+H���pxI��X{�����U%��!꣤87U�bń����DD��-zXlxV61EB     400     180>Y���E+�ݥFO-���ut9-Y��aܒ��`D�B�%�m����]�_Z�:	�>�+��<�Գ�[{r|xO�����1h�nZ����ъԿ�����N�~ʳ�"E| !�_�]�tA� 	�:Q� S��u�G.����m
|n�ҕ�Y��hP�E��0���+|�.*efaɼ8v��6��	��e5�b-h��c�YB�8J�p��â*�qY���*;��t��_k��Ł��_�����~�^`a~-H%0��@�ճH}<�*}Ҁ�~�K��x)��~��lbK��$B�f=5I �\o�ԩ�ѿ�Y�N+��� N�Ht�����`��尚T �[��Ǖ����4I��+��U�J������XlxV61EB     400      e0l3Jk��:6>�1�A�p^���=#*��<l����O+HfU�Տ���<X��l_��;�L�8��DC|{���v���H��]��)����k;v����О��zO4�E`ÁA�!�b�~1��2�<Ԍ�Vi�������ME-p��˨��� N�v}�2lOp��5�Mx��3`����eJ�~骣�4���:p��ǀ.c͸��"\�Ħ�L WMM[XlxV61EB     400      b0����4�&C����,X�s�Y�,���x���1�q�6ׯ�}I� �	�3�?<����(����0��V��2��9I�R����u��rc���V�ȁ�@@0��>֐��hDxЄ\�Z�n������t��6V�D�g�Pі�z2a��ò�4�T��،�Xw���qD�|ms��,�I�r��XlxV61EB     400     150��"| ܯ�lOGҧ&3�qj��{9��u1�W�ؕјe�hS�-ټ4����}�jȯ���`�ъ*.�o����������x&_Y���t}��#��Y���jC<05�\�?[&��]��}��}3�ֱI�ņ�Fo4��w�kf�ȫz�Owl_��쪦O攲C���=�U��J��m���H�Xz�v�?�*�����$V2}�0�!��t���~:�9�g�����c��Ô߽�C�I�_�������/���]�<�U�v0اD^}�I�<f��Y���F����|,�$��b��W���!����E�ڥ�r8�,�BV�����.�XlxV61EB     400      b0�҂u��7�Y�Uk�,�*�����dv��PUPZu{��qch$��hȕ�u��#'�+�+GA��do�'���Y;�O�=)��؉��J��T���+S��#ߺb��n���UN���HXC��>v�ԊZ}����]h�e��2�WZ+K���&���S�0Q��܏XlxV61EB     400     160'�h-�A!K����XG�N�����H.!���RaI���}`�="Ub�y &�z�e<�ku����	���F�x�Ŕ���f8$�%�HE;;����|���F;�����'���|o��UY�2&�W������X�?|��(��T�^)��Ы͟9{��u��#�d�}�Ĉ׽捛���{����GG��?m�jBѕ�K�g�2�u��#������
���F�*�!78§��3�ȶ�A����M�[��4j�vhdo ��ZAZ4�Y��q�*ݱ�V������
l'Ui��+���@��>96G��w�տ�!��C��_	��wQ��vw���:eXlxV61EB     400     140���e��3�eP�y�_ M�髍V������H�֢�������_�.\ ���S��� ��X���֥[�w>7ɏ�b��U8Y��J���][��6�[?���̍	Z!]2�Ex�K���jt(+�c($�(�R�mqXu�f3Z����2#�훻�|�;�r���Xڎ���c��@�7ޓ�����u�{�H���=9�a\}¡�ĞS����2ș�ѣ"H���򘷍G��?�'��W���V�
:�����������V#�#�s��G��A��:���fJX�1Q�Jw�	�`�Y@*�SZ�yٍ��7bԎXlxV61EB     400      b0�Bs���./��'@�ɼ��ő�E�lU���xc�RP�� ����='2t�h�8�Z�tb�B�²)m��D������F��h��XłD��'>~�Nt�f�ԝ�m�Dĺ"�jl�������8��s�?���,�=IA��B%��(
��� .���ym��Y�J�	;*���eXlxV61EB     400     180�4F�ZQvv���D���Z��s���[e��X3L�'�6����q<{F�pe��;�+C�c@�.=�9�1���!� žc�#:U��3�JՈi�%�n��a0�x��("Gj�����/�[�(4<�SGV�@��r�2!%����G��@�zPҶ���M��c�����K�կ��0�������X�U9S��6	�g���N��$%��V��f�E�蓌8c�n�7'i��:���O# �k�*yi�o�Λx�VсR%���%u,�x�,c���D��&�����N��a� ��_)����:��NG)>9�c."��Q,T�c�=Z�3xa��� tr*+����Z�:��Wz���U�	����"� �h�Hd���H������=�Q�XlxV61EB     400      b0G�/�𼢹����E�O���T��Bʜ�
��g8˸+Y�\�&7a 7_��IX!"�%���8V2�����>�U}�d��j�3��դ^��=@�/��[;�&:���:�$ڣ�Z�X]�Q��S%ozvu�3Ǟ�z�z� �D_�zO���ďK�5��>�{��iʔ�
i	BNhq��XlxV61EB     400      d0-	��-�]��x�T���e�I�?&��~j#�hpF=�d$�����%P�� ����V1R��'��P��dCD�������E�,r�ٴj
��͒6�׃V��K�o)	�q[��O�	-��S�~T�i}��!݌�"�Z���E�5��PFk �y/8\������l��OJ&���1��hR�ԝ)��x���*%�k��}eq0�,�
XlxV61EB     400     190�D<�!ȫ�� b E�߯����jC��\���sW���m��XO`�EO��;P��ĉYhv-~>�rR�A�@�M��D	��7��!���3�/�߀�
OPp��M�TH�0����T�/u2�1H`��/���jt��.p�]����=_��'U���W���;mR���{��nEG�oV!\�ٝ%��_�oG��>�t�5E���s"�	N}y!��s��W1�ȯ���3���LA�(%�h��
��(ё�4 �
���y�@������p��g�%kb$��;���<&��{���.J���M �^ښ�Y�>K��k�߉��\�ql��>��4�Y+&V�K٣��vƎ�Y���zueoߘn0�{pt{}��+���PXYp��N��fKXlxV61EB     400      b0�"L�����%�!]�/�8FFz�Y�����R]xc��U���
+���'�bM������9lR=��\� �3����(!ʐS
�o���"6NF߲���>4œ�0�p�+@�|�*�s%���)��xϸ��p!@u����/�6v��=��!>���ُ?m񬕺�T�XoXlxV61EB     400     140p�αEA���H<�B�B���A���x���b#K#��&(j5���y J�N���o瘺^"ՙ"���;��V}&�]�U2�䒰,R����[V[晼/�V��|F�2���8]>��?��(�n��l"��:~S%3���&j+T�G	0G�_�D��e�S@�X����s�%�2���^yH�R��Ga�\%
 �)�~g���S����[D?�:��R�G;�7"%ƫ�ܢ�o�I����sK�!^z1}W�hr��p�/�*�up=���-�o.BN��}�X.G����<�&k���,��%����eB����h��CXlxV61EB      10      20�k�.NO�'�aJ��Zt��g���ُ��zx