XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     170���Px�}�Y��}�iq*8��ǃN�DA��5�t�e�s�f���8�3�	1u9�ezs)���7���_�AW���bo������K�#�,���D�g跘�������A�9|2�kX�s��#�8�V]ƱjEiK�gR��R����j3��2�_����&�&�ǥ�Ɍ ��N��t��|��unӜ�0���S����gd3 ����������~2/E���4j�ך�NB�:�L����H��!�E�H��UC�O)<rF����i^f��OZpɛ)`���*h�����^F9�"�ߞ��"����׺��i����9��t�@�za,��9�@�2�H�9<_ԙm4�|cXlxV61EB     400     140`�Ȼ���^^8
0�o4�4��t� ��{�F˔"��$аpY���q���<>�kHU�Q�|DÛ����!�Դ�5շ�&N�ߴ�m����uFa���	�l�0BY�����֎�=�ȃ{�fY�y�yq{��v;JVB��/�� x �2B��}�ۥs�R��5\/;�?�[8k����J|7��j$7�n�8��,Hs����\.��C$橐߁�\�Ք4?��2/�L��d`�����Y7B�>g7h��/|�I����� <�]��{g�e�l��Q����wDI��I��H΃{��ڝ���M_�q�XlxV61EB     400     110�+�rY��e���(����@�o2?>��a���d��ӳ0+RX������VӪk������h��7}�����l����Ȟs@�A��r��Hw����Qq�:l)�,O4�H*�a�@eM��E��2r3H$�A��$�>\��5�5�R��=HDxol�GY�(�˨T����c���dz���y?�j���)�%��g2��Q��o�WT(��+����E�
����fOZ�h.=��lF�9�]��YТ�'��iD��Un�7i�ˑ�gY&nym[XlxV61EB     400     110![͗@:3q0�FFD�j�k-Ł+$ͮp��P���m[��`K�O��<>`R��� ���uS[(��Ĕ!~(h^`��-h�PR�e!���[�v,D��u�'9�����!�y(\8y���i��r/�2��w��������`��M����U�︭�T��Yº�z]��9@ts�V�&��q:4��3�=����".�)��c�T�2��!tF8+�MY�!�'��X�`A{X�U�.��U ��^I���������@����\#zh��+�t�XlxV61EB      9f      90R�$���޷b�y6�]�
op5*�]�w� y��{"���{Z�+��r�Iv躞���N}J�?�Gʇ�
���U]�xK�}����!����}|�F�2�p|�� CrB�	����VȨ.����ʫ�3��\